//*********************************************************************************************//
//    Project      : 16-Bit Multiplier Booth Recoder
//    File         : booth_recoder.v
//    Author       : Fasih-ud-Din Farrukh
//    Company      : Tsinghua University, Beijing, China
//    Start Date   : 
//    Last Updated : 
//    Version      : 0.1
//    Abstract     : This module implements ....
//
// 
//    Modification History:
//==============================================================================================
//    Date                       By                  Version                Change Description
//==============================================================================================
//    09th May, 2019           Rai Fasih              0.1                    Original Version
//*********************************************************************************************//

	`timescale 1ps/1ps                             

//------------------------------------------------------------------------------------------------------*/  
// Module of Booth recoder                                                                      
//------------------------------------------------------------------------------------------------------*/  

	module booth_recoder(//Inputs
											 recoderIn,
										 
		 									 //Outputs
											 recoderOut
											);

//------------------------------------------------------------------------------------------------------// 
// Input & Output Declarations                                                                  
//------------------------------------------------------------------------------------------------------// 
										
	input  [2:0] recoderIn;
	output [2:0] recoderOut;
	
//------------------------------------------------------------------------------------------------------// 
// Internal reg and wires declaration                                                                       
//------------------------------------------------------------------------------------------------------// 
	
	reg [2:0] recoderOut;

//------------------------------------------------------------------------------------------------------// 
// Case Statement                                                                  
//------------------------------------------------------------------------------------------------------//
	
	always @(recoderIn)
	begin
		case(recoderIn)
			3'b000: recoderOut = 3'b000; // 0
			3'b001: recoderOut = 3'b001; // 1
			3'b010: recoderOut = 3'b001; // 1
			3'b011: recoderOut = 3'b010; // 2
			3'b100: recoderOut = 3'b110; //-2
			3'b101: recoderOut = 3'b111; //-1
			3'b110: recoderOut = 3'b111; //-1
			3'b111: recoderOut = 3'b000; // 0
		 default: recoderOut = 3'bx;
		endcase
	end

//------------------------------------------------------------------------------------------------------// 
// End Module                                                                                      
//------------------------------------------------------------------------------------------------------// 
	
	endmodule										