VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO to_ALU_opt_TMR_KP_Voter
  CLASS BLOCK ;
  FOREIGN to_ALU_opt_TMR_KP_Voter ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.755 BY 261.475 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END CLK
  PIN COUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 200.640 250.755 201.240 ;
    END
  END COUT
  PIN DATA_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 257.475 55.110 261.475 ;
    END
  END DATA_IN
  PIN OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END OUT[0]
  PIN OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END OUT[10]
  PIN OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 257.475 193.570 261.475 ;
    END
  END OUT[11]
  PIN OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END OUT[12]
  PIN OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END OUT[13]
  PIN OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 142.840 250.755 143.440 ;
    END
  END OUT[14]
  PIN OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 257.475 248.310 261.475 ;
    END
  END OUT[15]
  PIN OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 257.475 138.830 261.475 ;
    END
  END OUT[1]
  PIN OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END OUT[2]
  PIN OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END OUT[3]
  PIN OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END OUT[4]
  PIN OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 173.440 250.755 174.040 ;
    END
  END OUT[5]
  PIN OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END OUT[6]
  PIN OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 54.440 250.755 55.040 ;
    END
  END OUT[7]
  PIN OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 257.475 167.810 261.475 ;
    END
  END OUT[8]
  PIN OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END OUT[9]
  PIN OUT_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 257.475 29.350 261.475 ;
    END
  END OUT_2[0]
  PIN OUT_2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END OUT_2[10]
  PIN OUT_2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 257.475 222.550 261.475 ;
    END
  END OUT_2[11]
  PIN OUT_2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 27.240 250.755 27.840 ;
    END
  END OUT_2[12]
  PIN OUT_2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END OUT_2[13]
  PIN OUT_2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END OUT_2[14]
  PIN OUT_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END OUT_2[1]
  PIN OUT_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 85.040 250.755 85.640 ;
    END
  END OUT_2[2]
  PIN OUT_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END OUT_2[3]
  PIN OUT_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END OUT_2[4]
  PIN OUT_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 231.240 250.755 231.840 ;
    END
  END OUT_2[5]
  PIN OUT_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 257.475 84.090 261.475 ;
    END
  END OUT_2[6]
  PIN OUT_2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 257.475 109.850 261.475 ;
    END
  END OUT_2[7]
  PIN OUT_2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END OUT_2[8]
  PIN OUT_2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END OUT_2[9]
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 257.475 0.370 261.475 ;
    END
  END RST
  PIN Ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.755 112.240 250.755 112.840 ;
    END
  END Ready
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 245.180 104.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 250.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 245.180 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 245.180 181.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 250.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 250.480 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 245.180 250.325 ;
      LAYER met1 ;
        RECT 0.070 10.640 248.330 250.480 ;
      LAYER met2 ;
        RECT 0.650 257.195 28.790 257.475 ;
        RECT 29.630 257.195 54.550 257.475 ;
        RECT 55.390 257.195 83.530 257.475 ;
        RECT 84.370 257.195 109.290 257.475 ;
        RECT 110.130 257.195 138.270 257.475 ;
        RECT 139.110 257.195 167.250 257.475 ;
        RECT 168.090 257.195 193.010 257.475 ;
        RECT 193.850 257.195 221.990 257.475 ;
        RECT 222.830 257.195 247.750 257.475 ;
        RECT 0.100 4.280 248.300 257.195 ;
        RECT 0.650 3.670 25.570 4.280 ;
        RECT 26.410 3.670 54.550 4.280 ;
        RECT 55.390 3.670 80.310 4.280 ;
        RECT 81.150 3.670 109.290 4.280 ;
        RECT 110.130 3.670 138.270 4.280 ;
        RECT 139.110 3.670 164.030 4.280 ;
        RECT 164.870 3.670 193.010 4.280 ;
        RECT 193.850 3.670 218.770 4.280 ;
        RECT 219.610 3.670 247.750 4.280 ;
      LAYER met3 ;
        RECT 4.000 232.240 246.755 250.405 ;
        RECT 4.400 230.840 246.355 232.240 ;
        RECT 4.000 205.040 246.755 230.840 ;
        RECT 4.400 203.640 246.755 205.040 ;
        RECT 4.000 201.640 246.755 203.640 ;
        RECT 4.000 200.240 246.355 201.640 ;
        RECT 4.000 174.440 246.755 200.240 ;
        RECT 4.400 173.040 246.355 174.440 ;
        RECT 4.000 147.240 246.755 173.040 ;
        RECT 4.400 145.840 246.755 147.240 ;
        RECT 4.000 143.840 246.755 145.840 ;
        RECT 4.000 142.440 246.355 143.840 ;
        RECT 4.000 116.640 246.755 142.440 ;
        RECT 4.400 115.240 246.755 116.640 ;
        RECT 4.000 113.240 246.755 115.240 ;
        RECT 4.000 111.840 246.355 113.240 ;
        RECT 4.000 86.040 246.755 111.840 ;
        RECT 4.400 84.640 246.355 86.040 ;
        RECT 4.000 58.840 246.755 84.640 ;
        RECT 4.400 57.440 246.755 58.840 ;
        RECT 4.000 55.440 246.755 57.440 ;
        RECT 4.000 54.040 246.355 55.440 ;
        RECT 4.000 28.240 246.755 54.040 ;
        RECT 4.400 26.840 246.355 28.240 ;
        RECT 4.000 10.715 246.755 26.840 ;
      LAYER met4 ;
        RECT 93.215 48.455 97.440 180.705 ;
        RECT 99.840 48.455 173.585 180.705 ;
  END
END to_ALU_opt_TMR_KP_Voter
END LIBRARY

