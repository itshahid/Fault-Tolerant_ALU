magic
tech sky130A
magscale 1 2
timestamp 1640855983
<< metal1 >>
rect 19518 700748 19524 700800
rect 19576 700788 19582 700800
rect 89162 700788 89168 700800
rect 19576 700760 89168 700788
rect 19576 700748 19582 700760
rect 89162 700748 89168 700760
rect 89220 700748 89226 700800
rect 76558 700680 76564 700732
rect 76616 700720 76622 700732
rect 154114 700720 154120 700732
rect 76616 700692 154120 700720
rect 76616 700680 76622 700692
rect 154114 700680 154120 700692
rect 154172 700680 154178 700732
rect 73798 700612 73804 700664
rect 73856 700652 73862 700664
rect 218974 700652 218980 700664
rect 73856 700624 218980 700652
rect 73856 700612 73862 700624
rect 218974 700612 218980 700624
rect 219032 700612 219038 700664
rect 17862 700544 17868 700596
rect 17920 700584 17926 700596
rect 283834 700584 283840 700596
rect 17920 700556 283840 700584
rect 17920 700544 17926 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 26142 700476 26148 700528
rect 26200 700516 26206 700528
rect 348786 700516 348792 700528
rect 26200 700488 348792 700516
rect 26200 700476 26206 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 70302 700408 70308 700460
rect 70360 700448 70366 700460
rect 413646 700448 413652 700460
rect 70360 700420 413652 700448
rect 70360 700408 70366 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 70026 700380 70032 700392
rect 24360 700352 70032 700380
rect 24360 700340 24366 700352
rect 70026 700340 70032 700352
rect 70084 700340 70090 700392
rect 72418 700340 72424 700392
rect 72476 700380 72482 700392
rect 478506 700380 478512 700392
rect 72476 700352 478512 700380
rect 72476 700340 72482 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 17770 700272 17776 700324
rect 17828 700312 17834 700324
rect 543458 700312 543464 700324
rect 17828 700284 543464 700312
rect 17828 700272 17834 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 17678 683136 17684 683188
rect 17736 683176 17742 683188
rect 580166 683176 580172 683188
rect 17736 683148 580172 683176
rect 17736 683136 17742 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 59262 630640 59268 630692
rect 59320 630680 59326 630692
rect 580166 630680 580172 630692
rect 59320 630652 580172 630680
rect 59320 630640 59326 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 2774 618400 2780 618452
rect 2832 618440 2838 618452
rect 6178 618440 6184 618452
rect 2832 618412 6184 618440
rect 2832 618400 2838 618412
rect 6178 618400 6184 618412
rect 6236 618400 6242 618452
rect 17586 524424 17592 524476
rect 17644 524464 17650 524476
rect 580166 524464 580172 524476
rect 17644 524436 580172 524464
rect 17644 524424 17650 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 7558 514808 7564 514820
rect 3384 514780 7564 514808
rect 3384 514768 3390 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 53742 470568 53748 470620
rect 53800 470608 53806 470620
rect 580166 470608 580172 470620
rect 53800 470580 580172 470608
rect 53800 470568 53806 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 72510 418140 72516 418192
rect 72568 418180 72574 418192
rect 580166 418180 580172 418192
rect 72568 418152 580172 418180
rect 72568 418140 72574 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 19426 364352 19432 364404
rect 19484 364392 19490 364404
rect 579614 364392 579620 364404
rect 19484 364364 579620 364392
rect 19484 364352 19490 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 2958 357416 2964 357468
rect 3016 357456 3022 357468
rect 69750 357456 69756 357468
rect 3016 357428 69756 357456
rect 3016 357416 3022 357428
rect 69750 357416 69756 357428
rect 69808 357416 69814 357468
rect 72602 311856 72608 311908
rect 72660 311896 72666 311908
rect 579982 311896 579988 311908
rect 72660 311868 579988 311896
rect 72660 311856 72666 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3050 304988 3056 305040
rect 3108 305028 3114 305040
rect 13078 305028 13084 305040
rect 3108 305000 13084 305028
rect 3108 304988 3114 305000
rect 13078 304988 13084 305000
rect 13136 304988 13142 305040
rect 17494 258068 17500 258120
rect 17552 258108 17558 258120
rect 580166 258108 580172 258120
rect 17552 258080 580172 258108
rect 17552 258068 17558 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3326 253920 3332 253972
rect 3384 253960 3390 253972
rect 15838 253960 15844 253972
rect 3384 253932 15844 253960
rect 3384 253920 3390 253932
rect 15838 253920 15844 253932
rect 15896 253920 15902 253972
rect 69842 218016 69848 218068
rect 69900 218056 69906 218068
rect 579890 218056 579896 218068
rect 69900 218028 579896 218056
rect 69900 218016 69906 218028
rect 579890 218016 579896 218028
rect 579948 218016 579954 218068
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 69934 201532 69940 201544
rect 3384 201504 69940 201532
rect 3384 201492 3390 201504
rect 69934 201492 69940 201504
rect 69992 201492 69998 201544
rect 17402 178032 17408 178084
rect 17460 178072 17466 178084
rect 580166 178072 580172 178084
rect 17460 178044 580172 178072
rect 17460 178032 17466 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 48222 137980 48228 138032
rect 48280 138020 48286 138032
rect 580166 138020 580172 138032
rect 48280 137992 580172 138020
rect 48280 137980 48286 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 83458 99356 83464 99408
rect 83516 99396 83522 99408
rect 580166 99396 580172 99408
rect 83516 99368 580172 99396
rect 83516 99356 83522 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 69658 75828 69664 75880
rect 69716 75868 69722 75880
rect 70302 75868 70308 75880
rect 69716 75840 70308 75868
rect 69716 75828 69722 75840
rect 70302 75828 70308 75840
rect 70360 75828 70366 75880
rect 3418 75284 3424 75336
rect 3476 75324 3482 75336
rect 36446 75324 36452 75336
rect 3476 75296 36452 75324
rect 3476 75284 3482 75296
rect 36446 75284 36452 75296
rect 36504 75284 36510 75336
rect 6178 75216 6184 75268
rect 6236 75256 6242 75268
rect 41598 75256 41604 75268
rect 6236 75228 41604 75256
rect 6236 75216 6242 75228
rect 41598 75216 41604 75228
rect 41656 75216 41662 75268
rect 3694 75148 3700 75200
rect 3752 75188 3758 75200
rect 64138 75188 64144 75200
rect 3752 75160 64144 75188
rect 3752 75148 3758 75160
rect 64138 75148 64144 75160
rect 64196 75148 64202 75200
rect 2682 74536 2688 74588
rect 2740 74576 2746 74588
rect 19702 74576 19708 74588
rect 2740 74548 19708 74576
rect 2740 74536 2746 74548
rect 19702 74536 19708 74548
rect 19760 74536 19766 74588
rect 72418 45568 72424 45620
rect 72476 45608 72482 45620
rect 579614 45608 579620 45620
rect 72476 45580 579620 45608
rect 72476 45568 72482 45580
rect 579614 45568 579620 45580
rect 579672 45568 579678 45620
rect 7558 44072 7564 44124
rect 7616 44112 7622 44124
rect 17770 44112 17776 44124
rect 7616 44084 17776 44112
rect 7616 44072 7622 44084
rect 17770 44072 17776 44084
rect 17828 44072 17834 44124
rect 71774 37068 71780 37120
rect 71832 37108 71838 37120
rect 73798 37108 73804 37120
rect 71832 37080 73804 37108
rect 71832 37068 71838 37080
rect 73798 37068 73804 37080
rect 73856 37068 73862 37120
rect 15838 17892 15844 17944
rect 15896 17932 15902 17944
rect 30650 17932 30656 17944
rect 15896 17904 30656 17932
rect 15896 17892 15902 17904
rect 30650 17892 30656 17904
rect 30708 17892 30714 17944
rect 36446 17892 36452 17944
rect 36504 17932 36510 17944
rect 580258 17932 580264 17944
rect 36504 17904 580264 17932
rect 36504 17892 36510 17904
rect 580258 17892 580264 17904
rect 580316 17892 580322 17944
rect 3602 17824 3608 17876
rect 3660 17864 3666 17876
rect 58342 17864 58348 17876
rect 3660 17836 58348 17864
rect 3660 17824 3666 17836
rect 58342 17824 58348 17836
rect 58400 17824 58406 17876
rect 64138 17824 64144 17876
rect 64196 17864 64202 17876
rect 64782 17864 64788 17876
rect 64196 17836 64788 17864
rect 64196 17824 64202 17836
rect 64782 17824 64788 17836
rect 64840 17824 64846 17876
rect 3510 17756 3516 17808
rect 3568 17796 3574 17808
rect 52546 17796 52552 17808
rect 3568 17768 52552 17796
rect 3568 17756 3574 17768
rect 52546 17756 52552 17768
rect 52604 17756 52610 17808
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 24854 17728 24860 17740
rect 13136 17700 24860 17728
rect 13136 17688 13142 17700
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 48038 17688 48044 17740
rect 48096 17728 48102 17740
rect 83458 17728 83464 17740
rect 48096 17700 83464 17728
rect 48096 17688 48102 17700
rect 83458 17688 83464 17700
rect 83516 17688 83522 17740
rect 42242 17620 42248 17672
rect 42300 17660 42306 17672
rect 76558 17660 76564 17672
rect 42300 17632 76564 17660
rect 42300 17620 42306 17632
rect 76558 17620 76564 17632
rect 76616 17620 76622 17672
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 64782 3408 64788 3460
rect 64840 3448 64846 3460
rect 579798 3448 579804 3460
rect 64840 3420 579804 3448
rect 64840 3408 64846 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
<< via1 >>
rect 19524 700748 19576 700800
rect 89168 700748 89220 700800
rect 76564 700680 76616 700732
rect 154120 700680 154172 700732
rect 73804 700612 73856 700664
rect 218980 700612 219032 700664
rect 17868 700544 17920 700596
rect 283840 700544 283892 700596
rect 26148 700476 26200 700528
rect 348792 700476 348844 700528
rect 70308 700408 70360 700460
rect 413652 700408 413704 700460
rect 24308 700340 24360 700392
rect 70032 700340 70084 700392
rect 72424 700340 72476 700392
rect 478512 700340 478564 700392
rect 17776 700272 17828 700324
rect 543464 700272 543516 700324
rect 17684 683136 17736 683188
rect 580172 683136 580224 683188
rect 59268 630640 59320 630692
rect 580172 630640 580224 630692
rect 2780 618400 2832 618452
rect 6184 618400 6236 618452
rect 17592 524424 17644 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 7564 514768 7616 514820
rect 53748 470568 53800 470620
rect 580172 470568 580224 470620
rect 72516 418140 72568 418192
rect 580172 418140 580224 418192
rect 19432 364352 19484 364404
rect 579620 364352 579672 364404
rect 2964 357416 3016 357468
rect 69756 357416 69808 357468
rect 72608 311856 72660 311908
rect 579988 311856 580040 311908
rect 3056 304988 3108 305040
rect 13084 304988 13136 305040
rect 17500 258068 17552 258120
rect 580172 258068 580224 258120
rect 3332 253920 3384 253972
rect 15844 253920 15896 253972
rect 69848 218016 69900 218068
rect 579896 218016 579948 218068
rect 3332 201492 3384 201544
rect 69940 201492 69992 201544
rect 17408 178032 17460 178084
rect 580172 178032 580224 178084
rect 48228 137980 48280 138032
rect 580172 137980 580224 138032
rect 83464 99356 83516 99408
rect 580172 99356 580224 99408
rect 69664 75828 69716 75880
rect 70308 75828 70360 75880
rect 3424 75284 3476 75336
rect 36452 75284 36504 75336
rect 6184 75216 6236 75268
rect 41604 75216 41656 75268
rect 3700 75148 3752 75200
rect 64144 75148 64196 75200
rect 2688 74536 2740 74588
rect 19708 74536 19760 74588
rect 72424 45568 72476 45620
rect 579620 45568 579672 45620
rect 7564 44072 7616 44124
rect 17776 44072 17828 44124
rect 71780 37068 71832 37120
rect 73804 37068 73856 37120
rect 15844 17892 15896 17944
rect 30656 17892 30708 17944
rect 36452 17892 36504 17944
rect 580264 17892 580316 17944
rect 3608 17824 3660 17876
rect 58348 17824 58400 17876
rect 64144 17824 64196 17876
rect 64788 17824 64840 17876
rect 3516 17756 3568 17808
rect 52552 17756 52604 17808
rect 13084 17688 13136 17740
rect 24860 17688 24912 17740
rect 48044 17688 48096 17740
rect 83464 17688 83516 17740
rect 42248 17620 42300 17672
rect 76564 17620 76616 17672
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 64788 3408 64840 3460
rect 579804 3408 579856 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 19524 700800 19576 700806
rect 19524 700742 19576 700748
rect 17868 700596 17920 700602
rect 17868 700538 17920 700544
rect 17776 700324 17828 700330
rect 17776 700266 17828 700272
rect 17684 683188 17736 683194
rect 17684 683130 17736 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2778 619168 2834 619177
rect 2778 619103 2834 619112
rect 2792 618458 2820 619103
rect 2780 618452 2832 618458
rect 2780 618394 2832 618400
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2962 358456 3018 358465
rect 2962 358391 3018 358400
rect 2976 357474 3004 358391
rect 2964 357468 3016 357474
rect 2964 357410 3016 357416
rect 3054 306232 3110 306241
rect 3054 306167 3110 306176
rect 3068 305046 3096 306167
rect 3056 305040 3108 305046
rect 3056 304982 3108 304988
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3344 253978 3372 254079
rect 3332 253972 3384 253978
rect 3332 253914 3384 253920
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3436 75342 3464 671191
rect 6184 618452 6236 618458
rect 6184 618394 6236 618400
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3424 75336 3476 75342
rect 3424 75278 3476 75284
rect 2688 74588 2740 74594
rect 2688 74530 2740 74536
rect 2700 3534 2728 74530
rect 3528 17814 3556 566879
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3620 17882 3648 462567
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 3712 75206 3740 410479
rect 6196 75274 6224 618394
rect 17592 524476 17644 524482
rect 17592 524418 17644 524424
rect 7564 514820 7616 514826
rect 7564 514762 7616 514768
rect 6184 75268 6236 75274
rect 6184 75210 6236 75216
rect 3700 75200 3752 75206
rect 3700 75142 3752 75148
rect 7576 44130 7604 514762
rect 13084 305040 13136 305046
rect 13084 304982 13136 304988
rect 7564 44124 7616 44130
rect 7564 44066 7616 44072
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 13096 17746 13124 304982
rect 17500 258120 17552 258126
rect 17500 258062 17552 258068
rect 15844 253972 15896 253978
rect 15844 253914 15896 253920
rect 15856 17950 15884 253914
rect 17408 178084 17460 178090
rect 17408 178026 17460 178032
rect 17420 66337 17448 178026
rect 17406 66328 17462 66337
rect 17406 66263 17462 66272
rect 17512 25537 17540 258062
rect 17604 54777 17632 524418
rect 17590 54768 17646 54777
rect 17590 54703 17646 54712
rect 17696 37097 17724 683130
rect 17788 49337 17816 700266
rect 17774 49328 17830 49337
rect 17774 49263 17830 49272
rect 17776 44124 17828 44130
rect 17776 44066 17828 44072
rect 17788 43217 17816 44066
rect 17774 43208 17830 43217
rect 17774 43143 17830 43152
rect 17682 37088 17738 37097
rect 17682 37023 17738 37032
rect 17880 31657 17908 700538
rect 19432 364404 19484 364410
rect 19432 364346 19484 364352
rect 19444 35894 19472 364346
rect 19536 60897 19564 700742
rect 24320 700398 24348 703520
rect 89180 700806 89208 703520
rect 89168 700800 89220 700806
rect 89168 700742 89220 700748
rect 154132 700738 154160 703520
rect 76564 700732 76616 700738
rect 76564 700674 76616 700680
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 73804 700664 73856 700670
rect 73804 700606 73856 700612
rect 26148 700528 26200 700534
rect 26148 700470 26200 700476
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 19708 74588 19760 74594
rect 19708 74530 19760 74536
rect 19720 72298 19748 74530
rect 26160 72298 26188 700470
rect 70308 700460 70360 700466
rect 70308 700402 70360 700408
rect 70032 700392 70084 700398
rect 70032 700334 70084 700340
rect 59268 630692 59320 630698
rect 59268 630634 59320 630640
rect 53748 470620 53800 470626
rect 53748 470562 53800 470568
rect 48228 138032 48280 138038
rect 48228 137974 48280 137980
rect 36452 75336 36504 75342
rect 36452 75278 36504 75284
rect 19720 72270 20056 72298
rect 25852 72270 26188 72298
rect 36464 72298 36492 75278
rect 41604 75268 41656 75274
rect 41604 75210 41656 75216
rect 41616 72298 41644 75210
rect 48240 74534 48268 137974
rect 48148 74506 48268 74534
rect 48148 72298 48176 74506
rect 53760 72298 53788 470562
rect 59280 74534 59308 630634
rect 69756 357468 69808 357474
rect 69756 357410 69808 357416
rect 69664 75880 69716 75886
rect 69664 75822 69716 75828
rect 64144 75200 64196 75206
rect 64144 75142 64196 75148
rect 59096 74506 59308 74534
rect 59096 72298 59124 74506
rect 36464 72270 36800 72298
rect 41616 72270 41952 72298
rect 47748 72270 48176 72298
rect 53544 72270 53788 72298
rect 58696 72270 59124 72298
rect 64156 72298 64184 75142
rect 69676 72298 69704 75822
rect 64156 72270 64492 72298
rect 69644 72270 69704 72298
rect 31298 71904 31354 71913
rect 31004 71862 31298 71890
rect 31298 71839 31354 71848
rect 19522 60888 19578 60897
rect 19522 60823 19578 60832
rect 19444 35866 19656 35894
rect 17866 31648 17922 31657
rect 17866 31583 17922 31592
rect 17498 25528 17554 25537
rect 17498 25463 17554 25472
rect 19628 20754 19656 35866
rect 69768 25945 69796 357410
rect 69848 218068 69900 218074
rect 69848 218010 69900 218016
rect 69754 25936 69810 25945
rect 69754 25871 69810 25880
rect 69860 20754 69888 218010
rect 69940 201544 69992 201550
rect 69940 201486 69992 201492
rect 69952 60625 69980 201486
rect 70044 66881 70072 700334
rect 70320 75886 70348 700402
rect 72424 700392 72476 700398
rect 72424 700334 72476 700340
rect 70308 75880 70360 75886
rect 70308 75822 70360 75828
rect 70030 66872 70086 66881
rect 70030 66807 70086 66816
rect 69938 60616 69994 60625
rect 69938 60551 69994 60560
rect 72436 48657 72464 700334
rect 72516 418192 72568 418198
rect 72516 418134 72568 418140
rect 72422 48648 72478 48657
rect 72422 48583 72478 48592
rect 72424 45620 72476 45626
rect 72424 45562 72476 45568
rect 72436 42537 72464 45562
rect 72422 42528 72478 42537
rect 72422 42463 72478 42472
rect 71780 37120 71832 37126
rect 71778 37088 71780 37097
rect 71832 37088 71834 37097
rect 71778 37023 71834 37032
rect 72528 30977 72556 418134
rect 72608 311908 72660 311914
rect 72608 311850 72660 311856
rect 72620 54777 72648 311850
rect 72606 54768 72662 54777
rect 72606 54703 72662 54712
rect 73816 37126 73844 700606
rect 73804 37120 73856 37126
rect 73804 37062 73856 37068
rect 72514 30968 72570 30977
rect 72514 30903 72570 30912
rect 19628 20726 20056 20754
rect 69644 20726 69888 20754
rect 24872 20046 25208 20074
rect 30668 20046 31004 20074
rect 36156 20046 36492 20074
rect 41952 20046 42288 20074
rect 47748 20046 48084 20074
rect 15844 17944 15896 17950
rect 15844 17886 15896 17892
rect 24872 17746 24900 20046
rect 30668 17950 30696 20046
rect 36464 17950 36492 20046
rect 30656 17944 30708 17950
rect 30656 17886 30708 17892
rect 36452 17944 36504 17950
rect 36452 17886 36504 17892
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 42260 17678 42288 20046
rect 48056 17746 48084 20046
rect 52564 20046 52900 20074
rect 58360 20046 58696 20074
rect 63848 20046 64184 20074
rect 52564 17814 52592 20046
rect 58360 17882 58388 20046
rect 64156 17882 64184 20046
rect 58348 17876 58400 17882
rect 58348 17818 58400 17824
rect 64144 17876 64196 17882
rect 64144 17818 64196 17824
rect 64788 17876 64840 17882
rect 64788 17818 64840 17824
rect 52552 17808 52604 17814
rect 52552 17750 52604 17756
rect 48044 17740 48096 17746
rect 48044 17682 48096 17688
rect 42248 17672 42300 17678
rect 42248 17614 42300 17620
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1688 480 1716 3470
rect 64800 3466 64828 17818
rect 76576 17678 76604 700674
rect 218992 700670 219020 703520
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 348804 700534 348832 703520
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 579908 218074 579936 218991
rect 579896 218068 579948 218074
rect 579896 218010 579948 218016
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 83464 99408 83516 99414
rect 83464 99350 83516 99356
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 83476 17746 83504 99350
rect 579618 46336 579674 46345
rect 579618 46271 579674 46280
rect 579632 45626 579660 46271
rect 579620 45620 579672 45626
rect 579620 45562 579672 45568
rect 580276 17950 580304 577623
rect 580264 17944 580316 17950
rect 580264 17886 580316 17892
rect 83464 17740 83516 17746
rect 83464 17682 83516 17688
rect 76564 17672 76616 17678
rect 76564 17614 76616 17620
rect 64788 3460 64840 3466
rect 64788 3402 64840 3408
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 671200 3478 671256
rect 2778 619112 2834 619168
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2962 358400 3018 358456
rect 3054 306176 3110 306232
rect 3330 254088 3386 254144
rect 3330 201864 3386 201920
rect 3514 566888 3570 566944
rect 3606 462576 3662 462632
rect 3698 410488 3754 410544
rect 17406 66272 17462 66328
rect 17590 54712 17646 54768
rect 17774 49272 17830 49328
rect 17774 43152 17830 43208
rect 17682 37032 17738 37088
rect 31298 71848 31354 71904
rect 19522 60832 19578 60888
rect 17866 31592 17922 31648
rect 17498 25472 17554 25528
rect 69754 25880 69810 25936
rect 70030 66816 70086 66872
rect 69938 60560 69994 60616
rect 72422 48592 72478 48648
rect 72422 42472 72478 42528
rect 71778 37068 71780 37088
rect 71780 37068 71832 37088
rect 71832 37068 71834 37088
rect 71778 37032 71834 37068
rect 72606 54712 72662 54768
rect 72514 30912 72570 30968
rect 580170 683848 580226 683904
rect 580170 630808 580226 630864
rect 580262 577632 580318 577688
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 471416 580226 471472
rect 580170 418240 580226 418296
rect 579618 365064 579674 365120
rect 579986 312024 580042 312080
rect 580170 258848 580226 258904
rect 579894 219000 579950 219056
rect 580170 179152 580226 179208
rect 580170 139304 580226 139360
rect 580170 99456 580226 99512
rect 579618 46280 579674 46336
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2957 358458 3023 358461
rect -960 358456 3023 358458
rect -960 358400 2962 358456
rect 3018 358400 3023 358456
rect -960 358398 3023 358400
rect -960 358308 480 358398
rect 2957 358395 3023 358398
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3049 306234 3115 306237
rect -960 306232 3115 306234
rect -960 306176 3054 306232
rect 3110 306176 3115 306232
rect -960 306174 3115 306176
rect -960 306084 480 306174
rect 3049 306171 3115 306174
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect 31293 71906 31359 71909
rect 31518 71906 31524 71908
rect 31293 71904 31524 71906
rect 31293 71848 31298 71904
rect 31354 71848 31524 71904
rect 31293 71846 31524 71848
rect 31293 71843 31359 71846
rect 31518 71844 31524 71846
rect 31588 71844 31594 71908
rect -960 71484 480 71724
rect 70025 66874 70091 66877
rect 69982 66872 70091 66874
rect 69982 66816 70030 66872
rect 70086 66816 70091 66872
rect 69982 66811 70091 66816
rect 17401 66330 17467 66333
rect 17401 66328 20148 66330
rect 17401 66272 17406 66328
rect 17462 66272 20148 66328
rect 69982 66300 70042 66811
rect 17401 66270 20148 66272
rect 17401 66267 17467 66270
rect 19517 60890 19583 60893
rect 19517 60888 20148 60890
rect 19517 60832 19522 60888
rect 19578 60832 20148 60888
rect 19517 60830 20148 60832
rect 19517 60827 19583 60830
rect 69933 60618 69999 60621
rect 69933 60616 70042 60618
rect 69933 60560 69938 60616
rect 69994 60560 70042 60616
rect 69933 60555 70042 60560
rect 69982 60180 70042 60555
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 17585 54770 17651 54773
rect 72601 54770 72667 54773
rect 17585 54768 20148 54770
rect 17585 54712 17590 54768
rect 17646 54712 20148 54768
rect 17585 54710 20148 54712
rect 70012 54768 72667 54770
rect 70012 54712 72606 54768
rect 72662 54712 72667 54768
rect 70012 54710 72667 54712
rect 17585 54707 17651 54710
rect 72601 54707 72667 54710
rect 17769 49330 17835 49333
rect 17769 49328 20148 49330
rect 17769 49272 17774 49328
rect 17830 49272 20148 49328
rect 17769 49270 20148 49272
rect 17769 49267 17835 49270
rect 72417 48650 72483 48653
rect 70012 48648 72483 48650
rect 70012 48592 72422 48648
rect 72478 48592 72483 48648
rect 70012 48590 72483 48592
rect 72417 48587 72483 48590
rect 579613 46338 579679 46341
rect 583520 46338 584960 46428
rect 579613 46336 584960 46338
rect 579613 46280 579618 46336
rect 579674 46280 584960 46336
rect 579613 46278 584960 46280
rect 579613 46275 579679 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 17769 43210 17835 43213
rect 17769 43208 20148 43210
rect 17769 43152 17774 43208
rect 17830 43152 20148 43208
rect 17769 43150 20148 43152
rect 17769 43147 17835 43150
rect 72417 42530 72483 42533
rect 70012 42528 72483 42530
rect 70012 42472 72422 42528
rect 72478 42472 72483 42528
rect 70012 42470 72483 42472
rect 72417 42467 72483 42470
rect 17677 37090 17743 37093
rect 71773 37090 71839 37093
rect 17677 37088 20148 37090
rect 17677 37032 17682 37088
rect 17738 37032 20148 37088
rect 17677 37030 20148 37032
rect 70012 37088 71839 37090
rect 70012 37032 71778 37088
rect 71834 37032 71839 37088
rect 70012 37030 71839 37032
rect 17677 37027 17743 37030
rect 71773 37027 71839 37030
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 17861 31650 17927 31653
rect 17861 31648 20148 31650
rect 17861 31592 17866 31648
rect 17922 31592 20148 31648
rect 17861 31590 20148 31592
rect 17861 31587 17927 31590
rect 72509 30970 72575 30973
rect 70012 30968 72575 30970
rect 70012 30912 72514 30968
rect 72570 30912 72575 30968
rect 70012 30910 72575 30912
rect 72509 30907 72575 30910
rect 69749 25938 69815 25941
rect 69749 25936 69858 25938
rect 69749 25880 69754 25936
rect 69810 25880 69858 25936
rect 69749 25875 69858 25880
rect 17493 25530 17559 25533
rect 17493 25528 20148 25530
rect 17493 25472 17498 25528
rect 17554 25472 20148 25528
rect 69798 25500 69858 25875
rect 17493 25470 20148 25472
rect 17493 25467 17559 25470
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 583520 6626 584960 6716
rect -960 6340 480 6580
rect 583342 6566 584960 6626
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect 31518 5612 31524 5676
rect 31588 5674 31594 5676
rect 583526 5674 583586 6430
rect 31588 5614 583586 5674
rect 31588 5612 31594 5614
<< via3 >>
rect 31524 71844 31588 71908
rect 31524 5612 31588 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 11954 710598 12574 711590
rect 11954 710362 11986 710598
rect 12222 710362 12306 710598
rect 12542 710362 12574 710598
rect 11954 710278 12574 710362
rect 11954 710042 11986 710278
rect 12222 710042 12306 710278
rect 12542 710042 12574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 8234 708678 8854 709670
rect 8234 708442 8266 708678
rect 8502 708442 8586 708678
rect 8822 708442 8854 708678
rect 8234 708358 8854 708442
rect 8234 708122 8266 708358
rect 8502 708122 8586 708358
rect 8822 708122 8854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 4514 706758 5134 707750
rect 4514 706522 4546 706758
rect 4782 706522 4866 706758
rect 5102 706522 5134 706758
rect 4514 706438 5134 706522
rect 4514 706202 4546 706438
rect 4782 706202 4866 706438
rect 5102 706202 5134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 794 704838 1414 705830
rect 794 704602 826 704838
rect 1062 704602 1146 704838
rect 1382 704602 1414 704838
rect 794 704518 1414 704602
rect 794 704282 826 704518
rect 1062 704282 1146 704518
rect 1382 704282 1414 704518
rect 794 687454 1414 704282
rect 794 687218 826 687454
rect 1062 687218 1146 687454
rect 1382 687218 1414 687454
rect 794 687134 1414 687218
rect 794 686898 826 687134
rect 1062 686898 1146 687134
rect 1382 686898 1414 687134
rect 794 651454 1414 686898
rect 794 651218 826 651454
rect 1062 651218 1146 651454
rect 1382 651218 1414 651454
rect 794 651134 1414 651218
rect 794 650898 826 651134
rect 1062 650898 1146 651134
rect 1382 650898 1414 651134
rect 794 615454 1414 650898
rect 794 615218 826 615454
rect 1062 615218 1146 615454
rect 1382 615218 1414 615454
rect 794 615134 1414 615218
rect 794 614898 826 615134
rect 1062 614898 1146 615134
rect 1382 614898 1414 615134
rect 794 579454 1414 614898
rect 794 579218 826 579454
rect 1062 579218 1146 579454
rect 1382 579218 1414 579454
rect 794 579134 1414 579218
rect 794 578898 826 579134
rect 1062 578898 1146 579134
rect 1382 578898 1414 579134
rect 794 543454 1414 578898
rect 794 543218 826 543454
rect 1062 543218 1146 543454
rect 1382 543218 1414 543454
rect 794 543134 1414 543218
rect 794 542898 826 543134
rect 1062 542898 1146 543134
rect 1382 542898 1414 543134
rect 794 507454 1414 542898
rect 794 507218 826 507454
rect 1062 507218 1146 507454
rect 1382 507218 1414 507454
rect 794 507134 1414 507218
rect 794 506898 826 507134
rect 1062 506898 1146 507134
rect 1382 506898 1414 507134
rect 794 471454 1414 506898
rect 794 471218 826 471454
rect 1062 471218 1146 471454
rect 1382 471218 1414 471454
rect 794 471134 1414 471218
rect 794 470898 826 471134
rect 1062 470898 1146 471134
rect 1382 470898 1414 471134
rect 794 435454 1414 470898
rect 794 435218 826 435454
rect 1062 435218 1146 435454
rect 1382 435218 1414 435454
rect 794 435134 1414 435218
rect 794 434898 826 435134
rect 1062 434898 1146 435134
rect 1382 434898 1414 435134
rect 794 399454 1414 434898
rect 794 399218 826 399454
rect 1062 399218 1146 399454
rect 1382 399218 1414 399454
rect 794 399134 1414 399218
rect 794 398898 826 399134
rect 1062 398898 1146 399134
rect 1382 398898 1414 399134
rect 794 363454 1414 398898
rect 794 363218 826 363454
rect 1062 363218 1146 363454
rect 1382 363218 1414 363454
rect 794 363134 1414 363218
rect 794 362898 826 363134
rect 1062 362898 1146 363134
rect 1382 362898 1414 363134
rect 794 327454 1414 362898
rect 794 327218 826 327454
rect 1062 327218 1146 327454
rect 1382 327218 1414 327454
rect 794 327134 1414 327218
rect 794 326898 826 327134
rect 1062 326898 1146 327134
rect 1382 326898 1414 327134
rect 794 291454 1414 326898
rect 794 291218 826 291454
rect 1062 291218 1146 291454
rect 1382 291218 1414 291454
rect 794 291134 1414 291218
rect 794 290898 826 291134
rect 1062 290898 1146 291134
rect 1382 290898 1414 291134
rect 794 255454 1414 290898
rect 794 255218 826 255454
rect 1062 255218 1146 255454
rect 1382 255218 1414 255454
rect 794 255134 1414 255218
rect 794 254898 826 255134
rect 1062 254898 1146 255134
rect 1382 254898 1414 255134
rect 794 219454 1414 254898
rect 794 219218 826 219454
rect 1062 219218 1146 219454
rect 1382 219218 1414 219454
rect 794 219134 1414 219218
rect 794 218898 826 219134
rect 1062 218898 1146 219134
rect 1382 218898 1414 219134
rect 794 183454 1414 218898
rect 794 183218 826 183454
rect 1062 183218 1146 183454
rect 1382 183218 1414 183454
rect 794 183134 1414 183218
rect 794 182898 826 183134
rect 1062 182898 1146 183134
rect 1382 182898 1414 183134
rect 794 147454 1414 182898
rect 794 147218 826 147454
rect 1062 147218 1146 147454
rect 1382 147218 1414 147454
rect 794 147134 1414 147218
rect 794 146898 826 147134
rect 1062 146898 1146 147134
rect 1382 146898 1414 147134
rect 794 111454 1414 146898
rect 794 111218 826 111454
rect 1062 111218 1146 111454
rect 1382 111218 1414 111454
rect 794 111134 1414 111218
rect 794 110898 826 111134
rect 1062 110898 1146 111134
rect 1382 110898 1414 111134
rect 794 75454 1414 110898
rect 794 75218 826 75454
rect 1062 75218 1146 75454
rect 1382 75218 1414 75454
rect 794 75134 1414 75218
rect 794 74898 826 75134
rect 1062 74898 1146 75134
rect 1382 74898 1414 75134
rect 794 39454 1414 74898
rect 794 39218 826 39454
rect 1062 39218 1146 39454
rect 1382 39218 1414 39454
rect 794 39134 1414 39218
rect 794 38898 826 39134
rect 1062 38898 1146 39134
rect 1382 38898 1414 39134
rect 794 3454 1414 38898
rect 794 3218 826 3454
rect 1062 3218 1146 3454
rect 1382 3218 1414 3454
rect 794 3134 1414 3218
rect 794 2898 826 3134
rect 1062 2898 1146 3134
rect 1382 2898 1414 3134
rect 794 -346 1414 2898
rect 794 -582 826 -346
rect 1062 -582 1146 -346
rect 1382 -582 1414 -346
rect 794 -666 1414 -582
rect 794 -902 826 -666
rect 1062 -902 1146 -666
rect 1382 -902 1414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 794 -1894 1414 -902
rect 4514 691174 5134 706202
rect 4514 690938 4546 691174
rect 4782 690938 4866 691174
rect 5102 690938 5134 691174
rect 4514 690854 5134 690938
rect 4514 690618 4546 690854
rect 4782 690618 4866 690854
rect 5102 690618 5134 690854
rect 4514 655174 5134 690618
rect 4514 654938 4546 655174
rect 4782 654938 4866 655174
rect 5102 654938 5134 655174
rect 4514 654854 5134 654938
rect 4514 654618 4546 654854
rect 4782 654618 4866 654854
rect 5102 654618 5134 654854
rect 4514 619174 5134 654618
rect 4514 618938 4546 619174
rect 4782 618938 4866 619174
rect 5102 618938 5134 619174
rect 4514 618854 5134 618938
rect 4514 618618 4546 618854
rect 4782 618618 4866 618854
rect 5102 618618 5134 618854
rect 4514 583174 5134 618618
rect 4514 582938 4546 583174
rect 4782 582938 4866 583174
rect 5102 582938 5134 583174
rect 4514 582854 5134 582938
rect 4514 582618 4546 582854
rect 4782 582618 4866 582854
rect 5102 582618 5134 582854
rect 4514 547174 5134 582618
rect 4514 546938 4546 547174
rect 4782 546938 4866 547174
rect 5102 546938 5134 547174
rect 4514 546854 5134 546938
rect 4514 546618 4546 546854
rect 4782 546618 4866 546854
rect 5102 546618 5134 546854
rect 4514 511174 5134 546618
rect 4514 510938 4546 511174
rect 4782 510938 4866 511174
rect 5102 510938 5134 511174
rect 4514 510854 5134 510938
rect 4514 510618 4546 510854
rect 4782 510618 4866 510854
rect 5102 510618 5134 510854
rect 4514 475174 5134 510618
rect 4514 474938 4546 475174
rect 4782 474938 4866 475174
rect 5102 474938 5134 475174
rect 4514 474854 5134 474938
rect 4514 474618 4546 474854
rect 4782 474618 4866 474854
rect 5102 474618 5134 474854
rect 4514 439174 5134 474618
rect 4514 438938 4546 439174
rect 4782 438938 4866 439174
rect 5102 438938 5134 439174
rect 4514 438854 5134 438938
rect 4514 438618 4546 438854
rect 4782 438618 4866 438854
rect 5102 438618 5134 438854
rect 4514 403174 5134 438618
rect 4514 402938 4546 403174
rect 4782 402938 4866 403174
rect 5102 402938 5134 403174
rect 4514 402854 5134 402938
rect 4514 402618 4546 402854
rect 4782 402618 4866 402854
rect 5102 402618 5134 402854
rect 4514 367174 5134 402618
rect 4514 366938 4546 367174
rect 4782 366938 4866 367174
rect 5102 366938 5134 367174
rect 4514 366854 5134 366938
rect 4514 366618 4546 366854
rect 4782 366618 4866 366854
rect 5102 366618 5134 366854
rect 4514 331174 5134 366618
rect 4514 330938 4546 331174
rect 4782 330938 4866 331174
rect 5102 330938 5134 331174
rect 4514 330854 5134 330938
rect 4514 330618 4546 330854
rect 4782 330618 4866 330854
rect 5102 330618 5134 330854
rect 4514 295174 5134 330618
rect 4514 294938 4546 295174
rect 4782 294938 4866 295174
rect 5102 294938 5134 295174
rect 4514 294854 5134 294938
rect 4514 294618 4546 294854
rect 4782 294618 4866 294854
rect 5102 294618 5134 294854
rect 4514 259174 5134 294618
rect 4514 258938 4546 259174
rect 4782 258938 4866 259174
rect 5102 258938 5134 259174
rect 4514 258854 5134 258938
rect 4514 258618 4546 258854
rect 4782 258618 4866 258854
rect 5102 258618 5134 258854
rect 4514 223174 5134 258618
rect 4514 222938 4546 223174
rect 4782 222938 4866 223174
rect 5102 222938 5134 223174
rect 4514 222854 5134 222938
rect 4514 222618 4546 222854
rect 4782 222618 4866 222854
rect 5102 222618 5134 222854
rect 4514 187174 5134 222618
rect 4514 186938 4546 187174
rect 4782 186938 4866 187174
rect 5102 186938 5134 187174
rect 4514 186854 5134 186938
rect 4514 186618 4546 186854
rect 4782 186618 4866 186854
rect 5102 186618 5134 186854
rect 4514 151174 5134 186618
rect 4514 150938 4546 151174
rect 4782 150938 4866 151174
rect 5102 150938 5134 151174
rect 4514 150854 5134 150938
rect 4514 150618 4546 150854
rect 4782 150618 4866 150854
rect 5102 150618 5134 150854
rect 4514 115174 5134 150618
rect 4514 114938 4546 115174
rect 4782 114938 4866 115174
rect 5102 114938 5134 115174
rect 4514 114854 5134 114938
rect 4514 114618 4546 114854
rect 4782 114618 4866 114854
rect 5102 114618 5134 114854
rect 4514 79174 5134 114618
rect 4514 78938 4546 79174
rect 4782 78938 4866 79174
rect 5102 78938 5134 79174
rect 4514 78854 5134 78938
rect 4514 78618 4546 78854
rect 4782 78618 4866 78854
rect 5102 78618 5134 78854
rect 4514 43174 5134 78618
rect 4514 42938 4546 43174
rect 4782 42938 4866 43174
rect 5102 42938 5134 43174
rect 4514 42854 5134 42938
rect 4514 42618 4546 42854
rect 4782 42618 4866 42854
rect 5102 42618 5134 42854
rect 4514 7174 5134 42618
rect 4514 6938 4546 7174
rect 4782 6938 4866 7174
rect 5102 6938 5134 7174
rect 4514 6854 5134 6938
rect 4514 6618 4546 6854
rect 4782 6618 4866 6854
rect 5102 6618 5134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 4514 -2266 5134 6618
rect 4514 -2502 4546 -2266
rect 4782 -2502 4866 -2266
rect 5102 -2502 5134 -2266
rect 4514 -2586 5134 -2502
rect 4514 -2822 4546 -2586
rect 4782 -2822 4866 -2586
rect 5102 -2822 5134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 4514 -3814 5134 -2822
rect 8234 694894 8854 708122
rect 8234 694658 8266 694894
rect 8502 694658 8586 694894
rect 8822 694658 8854 694894
rect 8234 694574 8854 694658
rect 8234 694338 8266 694574
rect 8502 694338 8586 694574
rect 8822 694338 8854 694574
rect 8234 658894 8854 694338
rect 8234 658658 8266 658894
rect 8502 658658 8586 658894
rect 8822 658658 8854 658894
rect 8234 658574 8854 658658
rect 8234 658338 8266 658574
rect 8502 658338 8586 658574
rect 8822 658338 8854 658574
rect 8234 622894 8854 658338
rect 8234 622658 8266 622894
rect 8502 622658 8586 622894
rect 8822 622658 8854 622894
rect 8234 622574 8854 622658
rect 8234 622338 8266 622574
rect 8502 622338 8586 622574
rect 8822 622338 8854 622574
rect 8234 586894 8854 622338
rect 8234 586658 8266 586894
rect 8502 586658 8586 586894
rect 8822 586658 8854 586894
rect 8234 586574 8854 586658
rect 8234 586338 8266 586574
rect 8502 586338 8586 586574
rect 8822 586338 8854 586574
rect 8234 550894 8854 586338
rect 8234 550658 8266 550894
rect 8502 550658 8586 550894
rect 8822 550658 8854 550894
rect 8234 550574 8854 550658
rect 8234 550338 8266 550574
rect 8502 550338 8586 550574
rect 8822 550338 8854 550574
rect 8234 514894 8854 550338
rect 8234 514658 8266 514894
rect 8502 514658 8586 514894
rect 8822 514658 8854 514894
rect 8234 514574 8854 514658
rect 8234 514338 8266 514574
rect 8502 514338 8586 514574
rect 8822 514338 8854 514574
rect 8234 478894 8854 514338
rect 8234 478658 8266 478894
rect 8502 478658 8586 478894
rect 8822 478658 8854 478894
rect 8234 478574 8854 478658
rect 8234 478338 8266 478574
rect 8502 478338 8586 478574
rect 8822 478338 8854 478574
rect 8234 442894 8854 478338
rect 8234 442658 8266 442894
rect 8502 442658 8586 442894
rect 8822 442658 8854 442894
rect 8234 442574 8854 442658
rect 8234 442338 8266 442574
rect 8502 442338 8586 442574
rect 8822 442338 8854 442574
rect 8234 406894 8854 442338
rect 8234 406658 8266 406894
rect 8502 406658 8586 406894
rect 8822 406658 8854 406894
rect 8234 406574 8854 406658
rect 8234 406338 8266 406574
rect 8502 406338 8586 406574
rect 8822 406338 8854 406574
rect 8234 370894 8854 406338
rect 8234 370658 8266 370894
rect 8502 370658 8586 370894
rect 8822 370658 8854 370894
rect 8234 370574 8854 370658
rect 8234 370338 8266 370574
rect 8502 370338 8586 370574
rect 8822 370338 8854 370574
rect 8234 334894 8854 370338
rect 8234 334658 8266 334894
rect 8502 334658 8586 334894
rect 8822 334658 8854 334894
rect 8234 334574 8854 334658
rect 8234 334338 8266 334574
rect 8502 334338 8586 334574
rect 8822 334338 8854 334574
rect 8234 298894 8854 334338
rect 8234 298658 8266 298894
rect 8502 298658 8586 298894
rect 8822 298658 8854 298894
rect 8234 298574 8854 298658
rect 8234 298338 8266 298574
rect 8502 298338 8586 298574
rect 8822 298338 8854 298574
rect 8234 262894 8854 298338
rect 8234 262658 8266 262894
rect 8502 262658 8586 262894
rect 8822 262658 8854 262894
rect 8234 262574 8854 262658
rect 8234 262338 8266 262574
rect 8502 262338 8586 262574
rect 8822 262338 8854 262574
rect 8234 226894 8854 262338
rect 8234 226658 8266 226894
rect 8502 226658 8586 226894
rect 8822 226658 8854 226894
rect 8234 226574 8854 226658
rect 8234 226338 8266 226574
rect 8502 226338 8586 226574
rect 8822 226338 8854 226574
rect 8234 190894 8854 226338
rect 8234 190658 8266 190894
rect 8502 190658 8586 190894
rect 8822 190658 8854 190894
rect 8234 190574 8854 190658
rect 8234 190338 8266 190574
rect 8502 190338 8586 190574
rect 8822 190338 8854 190574
rect 8234 154894 8854 190338
rect 8234 154658 8266 154894
rect 8502 154658 8586 154894
rect 8822 154658 8854 154894
rect 8234 154574 8854 154658
rect 8234 154338 8266 154574
rect 8502 154338 8586 154574
rect 8822 154338 8854 154574
rect 8234 118894 8854 154338
rect 8234 118658 8266 118894
rect 8502 118658 8586 118894
rect 8822 118658 8854 118894
rect 8234 118574 8854 118658
rect 8234 118338 8266 118574
rect 8502 118338 8586 118574
rect 8822 118338 8854 118574
rect 8234 82894 8854 118338
rect 8234 82658 8266 82894
rect 8502 82658 8586 82894
rect 8822 82658 8854 82894
rect 8234 82574 8854 82658
rect 8234 82338 8266 82574
rect 8502 82338 8586 82574
rect 8822 82338 8854 82574
rect 8234 46894 8854 82338
rect 8234 46658 8266 46894
rect 8502 46658 8586 46894
rect 8822 46658 8854 46894
rect 8234 46574 8854 46658
rect 8234 46338 8266 46574
rect 8502 46338 8586 46574
rect 8822 46338 8854 46574
rect 8234 10894 8854 46338
rect 8234 10658 8266 10894
rect 8502 10658 8586 10894
rect 8822 10658 8854 10894
rect 8234 10574 8854 10658
rect 8234 10338 8266 10574
rect 8502 10338 8586 10574
rect 8822 10338 8854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 8234 -4186 8854 10338
rect 10794 705798 11414 705830
rect 10794 705562 10826 705798
rect 11062 705562 11146 705798
rect 11382 705562 11414 705798
rect 10794 705478 11414 705562
rect 10794 705242 10826 705478
rect 11062 705242 11146 705478
rect 11382 705242 11414 705478
rect 10794 669454 11414 705242
rect 10794 669218 10826 669454
rect 11062 669218 11146 669454
rect 11382 669218 11414 669454
rect 10794 669134 11414 669218
rect 10794 668898 10826 669134
rect 11062 668898 11146 669134
rect 11382 668898 11414 669134
rect 10794 633454 11414 668898
rect 10794 633218 10826 633454
rect 11062 633218 11146 633454
rect 11382 633218 11414 633454
rect 10794 633134 11414 633218
rect 10794 632898 10826 633134
rect 11062 632898 11146 633134
rect 11382 632898 11414 633134
rect 10794 597454 11414 632898
rect 10794 597218 10826 597454
rect 11062 597218 11146 597454
rect 11382 597218 11414 597454
rect 10794 597134 11414 597218
rect 10794 596898 10826 597134
rect 11062 596898 11146 597134
rect 11382 596898 11414 597134
rect 10794 561454 11414 596898
rect 10794 561218 10826 561454
rect 11062 561218 11146 561454
rect 11382 561218 11414 561454
rect 10794 561134 11414 561218
rect 10794 560898 10826 561134
rect 11062 560898 11146 561134
rect 11382 560898 11414 561134
rect 10794 525454 11414 560898
rect 10794 525218 10826 525454
rect 11062 525218 11146 525454
rect 11382 525218 11414 525454
rect 10794 525134 11414 525218
rect 10794 524898 10826 525134
rect 11062 524898 11146 525134
rect 11382 524898 11414 525134
rect 10794 489454 11414 524898
rect 10794 489218 10826 489454
rect 11062 489218 11146 489454
rect 11382 489218 11414 489454
rect 10794 489134 11414 489218
rect 10794 488898 10826 489134
rect 11062 488898 11146 489134
rect 11382 488898 11414 489134
rect 10794 453454 11414 488898
rect 10794 453218 10826 453454
rect 11062 453218 11146 453454
rect 11382 453218 11414 453454
rect 10794 453134 11414 453218
rect 10794 452898 10826 453134
rect 11062 452898 11146 453134
rect 11382 452898 11414 453134
rect 10794 417454 11414 452898
rect 10794 417218 10826 417454
rect 11062 417218 11146 417454
rect 11382 417218 11414 417454
rect 10794 417134 11414 417218
rect 10794 416898 10826 417134
rect 11062 416898 11146 417134
rect 11382 416898 11414 417134
rect 10794 381454 11414 416898
rect 10794 381218 10826 381454
rect 11062 381218 11146 381454
rect 11382 381218 11414 381454
rect 10794 381134 11414 381218
rect 10794 380898 10826 381134
rect 11062 380898 11146 381134
rect 11382 380898 11414 381134
rect 10794 345454 11414 380898
rect 10794 345218 10826 345454
rect 11062 345218 11146 345454
rect 11382 345218 11414 345454
rect 10794 345134 11414 345218
rect 10794 344898 10826 345134
rect 11062 344898 11146 345134
rect 11382 344898 11414 345134
rect 10794 309454 11414 344898
rect 10794 309218 10826 309454
rect 11062 309218 11146 309454
rect 11382 309218 11414 309454
rect 10794 309134 11414 309218
rect 10794 308898 10826 309134
rect 11062 308898 11146 309134
rect 11382 308898 11414 309134
rect 10794 273454 11414 308898
rect 10794 273218 10826 273454
rect 11062 273218 11146 273454
rect 11382 273218 11414 273454
rect 10794 273134 11414 273218
rect 10794 272898 10826 273134
rect 11062 272898 11146 273134
rect 11382 272898 11414 273134
rect 10794 237454 11414 272898
rect 10794 237218 10826 237454
rect 11062 237218 11146 237454
rect 11382 237218 11414 237454
rect 10794 237134 11414 237218
rect 10794 236898 10826 237134
rect 11062 236898 11146 237134
rect 11382 236898 11414 237134
rect 10794 201454 11414 236898
rect 10794 201218 10826 201454
rect 11062 201218 11146 201454
rect 11382 201218 11414 201454
rect 10794 201134 11414 201218
rect 10794 200898 10826 201134
rect 11062 200898 11146 201134
rect 11382 200898 11414 201134
rect 10794 165454 11414 200898
rect 10794 165218 10826 165454
rect 11062 165218 11146 165454
rect 11382 165218 11414 165454
rect 10794 165134 11414 165218
rect 10794 164898 10826 165134
rect 11062 164898 11146 165134
rect 11382 164898 11414 165134
rect 10794 129454 11414 164898
rect 10794 129218 10826 129454
rect 11062 129218 11146 129454
rect 11382 129218 11414 129454
rect 10794 129134 11414 129218
rect 10794 128898 10826 129134
rect 11062 128898 11146 129134
rect 11382 128898 11414 129134
rect 10794 93454 11414 128898
rect 10794 93218 10826 93454
rect 11062 93218 11146 93454
rect 11382 93218 11414 93454
rect 10794 93134 11414 93218
rect 10794 92898 10826 93134
rect 11062 92898 11146 93134
rect 11382 92898 11414 93134
rect 10794 57454 11414 92898
rect 10794 57218 10826 57454
rect 11062 57218 11146 57454
rect 11382 57218 11414 57454
rect 10794 57134 11414 57218
rect 10794 56898 10826 57134
rect 11062 56898 11146 57134
rect 11382 56898 11414 57134
rect 10794 21454 11414 56898
rect 10794 21218 10826 21454
rect 11062 21218 11146 21454
rect 11382 21218 11414 21454
rect 10794 21134 11414 21218
rect 10794 20898 10826 21134
rect 11062 20898 11146 21134
rect 11382 20898 11414 21134
rect 10794 -1306 11414 20898
rect 10794 -1542 10826 -1306
rect 11062 -1542 11146 -1306
rect 11382 -1542 11414 -1306
rect 10794 -1626 11414 -1542
rect 10794 -1862 10826 -1626
rect 11062 -1862 11146 -1626
rect 11382 -1862 11414 -1626
rect 10794 -1894 11414 -1862
rect 11954 698614 12574 710042
rect 21954 711558 22574 711590
rect 21954 711322 21986 711558
rect 22222 711322 22306 711558
rect 22542 711322 22574 711558
rect 21954 711238 22574 711322
rect 21954 711002 21986 711238
rect 22222 711002 22306 711238
rect 22542 711002 22574 711238
rect 18234 709638 18854 709670
rect 18234 709402 18266 709638
rect 18502 709402 18586 709638
rect 18822 709402 18854 709638
rect 18234 709318 18854 709402
rect 18234 709082 18266 709318
rect 18502 709082 18586 709318
rect 18822 709082 18854 709318
rect 11954 698378 11986 698614
rect 12222 698378 12306 698614
rect 12542 698378 12574 698614
rect 11954 698294 12574 698378
rect 11954 698058 11986 698294
rect 12222 698058 12306 698294
rect 12542 698058 12574 698294
rect 11954 662614 12574 698058
rect 11954 662378 11986 662614
rect 12222 662378 12306 662614
rect 12542 662378 12574 662614
rect 11954 662294 12574 662378
rect 11954 662058 11986 662294
rect 12222 662058 12306 662294
rect 12542 662058 12574 662294
rect 11954 626614 12574 662058
rect 11954 626378 11986 626614
rect 12222 626378 12306 626614
rect 12542 626378 12574 626614
rect 11954 626294 12574 626378
rect 11954 626058 11986 626294
rect 12222 626058 12306 626294
rect 12542 626058 12574 626294
rect 11954 590614 12574 626058
rect 11954 590378 11986 590614
rect 12222 590378 12306 590614
rect 12542 590378 12574 590614
rect 11954 590294 12574 590378
rect 11954 590058 11986 590294
rect 12222 590058 12306 590294
rect 12542 590058 12574 590294
rect 11954 554614 12574 590058
rect 11954 554378 11986 554614
rect 12222 554378 12306 554614
rect 12542 554378 12574 554614
rect 11954 554294 12574 554378
rect 11954 554058 11986 554294
rect 12222 554058 12306 554294
rect 12542 554058 12574 554294
rect 11954 518614 12574 554058
rect 11954 518378 11986 518614
rect 12222 518378 12306 518614
rect 12542 518378 12574 518614
rect 11954 518294 12574 518378
rect 11954 518058 11986 518294
rect 12222 518058 12306 518294
rect 12542 518058 12574 518294
rect 11954 482614 12574 518058
rect 11954 482378 11986 482614
rect 12222 482378 12306 482614
rect 12542 482378 12574 482614
rect 11954 482294 12574 482378
rect 11954 482058 11986 482294
rect 12222 482058 12306 482294
rect 12542 482058 12574 482294
rect 11954 446614 12574 482058
rect 11954 446378 11986 446614
rect 12222 446378 12306 446614
rect 12542 446378 12574 446614
rect 11954 446294 12574 446378
rect 11954 446058 11986 446294
rect 12222 446058 12306 446294
rect 12542 446058 12574 446294
rect 11954 410614 12574 446058
rect 11954 410378 11986 410614
rect 12222 410378 12306 410614
rect 12542 410378 12574 410614
rect 11954 410294 12574 410378
rect 11954 410058 11986 410294
rect 12222 410058 12306 410294
rect 12542 410058 12574 410294
rect 11954 374614 12574 410058
rect 11954 374378 11986 374614
rect 12222 374378 12306 374614
rect 12542 374378 12574 374614
rect 11954 374294 12574 374378
rect 11954 374058 11986 374294
rect 12222 374058 12306 374294
rect 12542 374058 12574 374294
rect 11954 338614 12574 374058
rect 11954 338378 11986 338614
rect 12222 338378 12306 338614
rect 12542 338378 12574 338614
rect 11954 338294 12574 338378
rect 11954 338058 11986 338294
rect 12222 338058 12306 338294
rect 12542 338058 12574 338294
rect 11954 302614 12574 338058
rect 11954 302378 11986 302614
rect 12222 302378 12306 302614
rect 12542 302378 12574 302614
rect 11954 302294 12574 302378
rect 11954 302058 11986 302294
rect 12222 302058 12306 302294
rect 12542 302058 12574 302294
rect 11954 266614 12574 302058
rect 11954 266378 11986 266614
rect 12222 266378 12306 266614
rect 12542 266378 12574 266614
rect 11954 266294 12574 266378
rect 11954 266058 11986 266294
rect 12222 266058 12306 266294
rect 12542 266058 12574 266294
rect 11954 230614 12574 266058
rect 11954 230378 11986 230614
rect 12222 230378 12306 230614
rect 12542 230378 12574 230614
rect 11954 230294 12574 230378
rect 11954 230058 11986 230294
rect 12222 230058 12306 230294
rect 12542 230058 12574 230294
rect 11954 194614 12574 230058
rect 11954 194378 11986 194614
rect 12222 194378 12306 194614
rect 12542 194378 12574 194614
rect 11954 194294 12574 194378
rect 11954 194058 11986 194294
rect 12222 194058 12306 194294
rect 12542 194058 12574 194294
rect 11954 158614 12574 194058
rect 11954 158378 11986 158614
rect 12222 158378 12306 158614
rect 12542 158378 12574 158614
rect 11954 158294 12574 158378
rect 11954 158058 11986 158294
rect 12222 158058 12306 158294
rect 12542 158058 12574 158294
rect 11954 122614 12574 158058
rect 11954 122378 11986 122614
rect 12222 122378 12306 122614
rect 12542 122378 12574 122614
rect 11954 122294 12574 122378
rect 11954 122058 11986 122294
rect 12222 122058 12306 122294
rect 12542 122058 12574 122294
rect 11954 86614 12574 122058
rect 11954 86378 11986 86614
rect 12222 86378 12306 86614
rect 12542 86378 12574 86614
rect 11954 86294 12574 86378
rect 11954 86058 11986 86294
rect 12222 86058 12306 86294
rect 12542 86058 12574 86294
rect 11954 50614 12574 86058
rect 11954 50378 11986 50614
rect 12222 50378 12306 50614
rect 12542 50378 12574 50614
rect 11954 50294 12574 50378
rect 11954 50058 11986 50294
rect 12222 50058 12306 50294
rect 12542 50058 12574 50294
rect 11954 14614 12574 50058
rect 11954 14378 11986 14614
rect 12222 14378 12306 14614
rect 12542 14378 12574 14614
rect 11954 14294 12574 14378
rect 11954 14058 11986 14294
rect 12222 14058 12306 14294
rect 12542 14058 12574 14294
rect 8234 -4422 8266 -4186
rect 8502 -4422 8586 -4186
rect 8822 -4422 8854 -4186
rect 8234 -4506 8854 -4422
rect 8234 -4742 8266 -4506
rect 8502 -4742 8586 -4506
rect 8822 -4742 8854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 8234 -5734 8854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 11954 -6106 12574 14058
rect 14514 707718 15134 707750
rect 14514 707482 14546 707718
rect 14782 707482 14866 707718
rect 15102 707482 15134 707718
rect 14514 707398 15134 707482
rect 14514 707162 14546 707398
rect 14782 707162 14866 707398
rect 15102 707162 15134 707398
rect 14514 673174 15134 707162
rect 14514 672938 14546 673174
rect 14782 672938 14866 673174
rect 15102 672938 15134 673174
rect 14514 672854 15134 672938
rect 14514 672618 14546 672854
rect 14782 672618 14866 672854
rect 15102 672618 15134 672854
rect 14514 637174 15134 672618
rect 14514 636938 14546 637174
rect 14782 636938 14866 637174
rect 15102 636938 15134 637174
rect 14514 636854 15134 636938
rect 14514 636618 14546 636854
rect 14782 636618 14866 636854
rect 15102 636618 15134 636854
rect 14514 601174 15134 636618
rect 14514 600938 14546 601174
rect 14782 600938 14866 601174
rect 15102 600938 15134 601174
rect 14514 600854 15134 600938
rect 14514 600618 14546 600854
rect 14782 600618 14866 600854
rect 15102 600618 15134 600854
rect 14514 565174 15134 600618
rect 14514 564938 14546 565174
rect 14782 564938 14866 565174
rect 15102 564938 15134 565174
rect 14514 564854 15134 564938
rect 14514 564618 14546 564854
rect 14782 564618 14866 564854
rect 15102 564618 15134 564854
rect 14514 529174 15134 564618
rect 14514 528938 14546 529174
rect 14782 528938 14866 529174
rect 15102 528938 15134 529174
rect 14514 528854 15134 528938
rect 14514 528618 14546 528854
rect 14782 528618 14866 528854
rect 15102 528618 15134 528854
rect 14514 493174 15134 528618
rect 14514 492938 14546 493174
rect 14782 492938 14866 493174
rect 15102 492938 15134 493174
rect 14514 492854 15134 492938
rect 14514 492618 14546 492854
rect 14782 492618 14866 492854
rect 15102 492618 15134 492854
rect 14514 457174 15134 492618
rect 14514 456938 14546 457174
rect 14782 456938 14866 457174
rect 15102 456938 15134 457174
rect 14514 456854 15134 456938
rect 14514 456618 14546 456854
rect 14782 456618 14866 456854
rect 15102 456618 15134 456854
rect 14514 421174 15134 456618
rect 14514 420938 14546 421174
rect 14782 420938 14866 421174
rect 15102 420938 15134 421174
rect 14514 420854 15134 420938
rect 14514 420618 14546 420854
rect 14782 420618 14866 420854
rect 15102 420618 15134 420854
rect 14514 385174 15134 420618
rect 14514 384938 14546 385174
rect 14782 384938 14866 385174
rect 15102 384938 15134 385174
rect 14514 384854 15134 384938
rect 14514 384618 14546 384854
rect 14782 384618 14866 384854
rect 15102 384618 15134 384854
rect 14514 349174 15134 384618
rect 14514 348938 14546 349174
rect 14782 348938 14866 349174
rect 15102 348938 15134 349174
rect 14514 348854 15134 348938
rect 14514 348618 14546 348854
rect 14782 348618 14866 348854
rect 15102 348618 15134 348854
rect 14514 313174 15134 348618
rect 14514 312938 14546 313174
rect 14782 312938 14866 313174
rect 15102 312938 15134 313174
rect 14514 312854 15134 312938
rect 14514 312618 14546 312854
rect 14782 312618 14866 312854
rect 15102 312618 15134 312854
rect 14514 277174 15134 312618
rect 14514 276938 14546 277174
rect 14782 276938 14866 277174
rect 15102 276938 15134 277174
rect 14514 276854 15134 276938
rect 14514 276618 14546 276854
rect 14782 276618 14866 276854
rect 15102 276618 15134 276854
rect 14514 241174 15134 276618
rect 14514 240938 14546 241174
rect 14782 240938 14866 241174
rect 15102 240938 15134 241174
rect 14514 240854 15134 240938
rect 14514 240618 14546 240854
rect 14782 240618 14866 240854
rect 15102 240618 15134 240854
rect 14514 205174 15134 240618
rect 14514 204938 14546 205174
rect 14782 204938 14866 205174
rect 15102 204938 15134 205174
rect 14514 204854 15134 204938
rect 14514 204618 14546 204854
rect 14782 204618 14866 204854
rect 15102 204618 15134 204854
rect 14514 169174 15134 204618
rect 14514 168938 14546 169174
rect 14782 168938 14866 169174
rect 15102 168938 15134 169174
rect 14514 168854 15134 168938
rect 14514 168618 14546 168854
rect 14782 168618 14866 168854
rect 15102 168618 15134 168854
rect 14514 133174 15134 168618
rect 14514 132938 14546 133174
rect 14782 132938 14866 133174
rect 15102 132938 15134 133174
rect 14514 132854 15134 132938
rect 14514 132618 14546 132854
rect 14782 132618 14866 132854
rect 15102 132618 15134 132854
rect 14514 97174 15134 132618
rect 14514 96938 14546 97174
rect 14782 96938 14866 97174
rect 15102 96938 15134 97174
rect 14514 96854 15134 96938
rect 14514 96618 14546 96854
rect 14782 96618 14866 96854
rect 15102 96618 15134 96854
rect 14514 61174 15134 96618
rect 18234 676894 18854 709082
rect 18234 676658 18266 676894
rect 18502 676658 18586 676894
rect 18822 676658 18854 676894
rect 18234 676574 18854 676658
rect 18234 676338 18266 676574
rect 18502 676338 18586 676574
rect 18822 676338 18854 676574
rect 18234 640894 18854 676338
rect 18234 640658 18266 640894
rect 18502 640658 18586 640894
rect 18822 640658 18854 640894
rect 18234 640574 18854 640658
rect 18234 640338 18266 640574
rect 18502 640338 18586 640574
rect 18822 640338 18854 640574
rect 18234 604894 18854 640338
rect 18234 604658 18266 604894
rect 18502 604658 18586 604894
rect 18822 604658 18854 604894
rect 18234 604574 18854 604658
rect 18234 604338 18266 604574
rect 18502 604338 18586 604574
rect 18822 604338 18854 604574
rect 18234 568894 18854 604338
rect 18234 568658 18266 568894
rect 18502 568658 18586 568894
rect 18822 568658 18854 568894
rect 18234 568574 18854 568658
rect 18234 568338 18266 568574
rect 18502 568338 18586 568574
rect 18822 568338 18854 568574
rect 18234 532894 18854 568338
rect 18234 532658 18266 532894
rect 18502 532658 18586 532894
rect 18822 532658 18854 532894
rect 18234 532574 18854 532658
rect 18234 532338 18266 532574
rect 18502 532338 18586 532574
rect 18822 532338 18854 532574
rect 18234 496894 18854 532338
rect 18234 496658 18266 496894
rect 18502 496658 18586 496894
rect 18822 496658 18854 496894
rect 18234 496574 18854 496658
rect 18234 496338 18266 496574
rect 18502 496338 18586 496574
rect 18822 496338 18854 496574
rect 18234 460894 18854 496338
rect 18234 460658 18266 460894
rect 18502 460658 18586 460894
rect 18822 460658 18854 460894
rect 18234 460574 18854 460658
rect 18234 460338 18266 460574
rect 18502 460338 18586 460574
rect 18822 460338 18854 460574
rect 18234 424894 18854 460338
rect 18234 424658 18266 424894
rect 18502 424658 18586 424894
rect 18822 424658 18854 424894
rect 18234 424574 18854 424658
rect 18234 424338 18266 424574
rect 18502 424338 18586 424574
rect 18822 424338 18854 424574
rect 18234 388894 18854 424338
rect 18234 388658 18266 388894
rect 18502 388658 18586 388894
rect 18822 388658 18854 388894
rect 18234 388574 18854 388658
rect 18234 388338 18266 388574
rect 18502 388338 18586 388574
rect 18822 388338 18854 388574
rect 18234 352894 18854 388338
rect 18234 352658 18266 352894
rect 18502 352658 18586 352894
rect 18822 352658 18854 352894
rect 18234 352574 18854 352658
rect 18234 352338 18266 352574
rect 18502 352338 18586 352574
rect 18822 352338 18854 352574
rect 18234 316894 18854 352338
rect 18234 316658 18266 316894
rect 18502 316658 18586 316894
rect 18822 316658 18854 316894
rect 18234 316574 18854 316658
rect 18234 316338 18266 316574
rect 18502 316338 18586 316574
rect 18822 316338 18854 316574
rect 18234 280894 18854 316338
rect 18234 280658 18266 280894
rect 18502 280658 18586 280894
rect 18822 280658 18854 280894
rect 18234 280574 18854 280658
rect 18234 280338 18266 280574
rect 18502 280338 18586 280574
rect 18822 280338 18854 280574
rect 18234 244894 18854 280338
rect 18234 244658 18266 244894
rect 18502 244658 18586 244894
rect 18822 244658 18854 244894
rect 18234 244574 18854 244658
rect 18234 244338 18266 244574
rect 18502 244338 18586 244574
rect 18822 244338 18854 244574
rect 18234 208894 18854 244338
rect 18234 208658 18266 208894
rect 18502 208658 18586 208894
rect 18822 208658 18854 208894
rect 18234 208574 18854 208658
rect 18234 208338 18266 208574
rect 18502 208338 18586 208574
rect 18822 208338 18854 208574
rect 18234 172894 18854 208338
rect 18234 172658 18266 172894
rect 18502 172658 18586 172894
rect 18822 172658 18854 172894
rect 18234 172574 18854 172658
rect 18234 172338 18266 172574
rect 18502 172338 18586 172574
rect 18822 172338 18854 172574
rect 18234 136894 18854 172338
rect 18234 136658 18266 136894
rect 18502 136658 18586 136894
rect 18822 136658 18854 136894
rect 18234 136574 18854 136658
rect 18234 136338 18266 136574
rect 18502 136338 18586 136574
rect 18822 136338 18854 136574
rect 18234 100894 18854 136338
rect 18234 100658 18266 100894
rect 18502 100658 18586 100894
rect 18822 100658 18854 100894
rect 18234 100574 18854 100658
rect 18234 100338 18266 100574
rect 18502 100338 18586 100574
rect 18822 100338 18854 100574
rect 18234 74295 18854 100338
rect 20794 704838 21414 705830
rect 20794 704602 20826 704838
rect 21062 704602 21146 704838
rect 21382 704602 21414 704838
rect 20794 704518 21414 704602
rect 20794 704282 20826 704518
rect 21062 704282 21146 704518
rect 21382 704282 21414 704518
rect 20794 687454 21414 704282
rect 20794 687218 20826 687454
rect 21062 687218 21146 687454
rect 21382 687218 21414 687454
rect 20794 687134 21414 687218
rect 20794 686898 20826 687134
rect 21062 686898 21146 687134
rect 21382 686898 21414 687134
rect 20794 651454 21414 686898
rect 20794 651218 20826 651454
rect 21062 651218 21146 651454
rect 21382 651218 21414 651454
rect 20794 651134 21414 651218
rect 20794 650898 20826 651134
rect 21062 650898 21146 651134
rect 21382 650898 21414 651134
rect 20794 615454 21414 650898
rect 20794 615218 20826 615454
rect 21062 615218 21146 615454
rect 21382 615218 21414 615454
rect 20794 615134 21414 615218
rect 20794 614898 20826 615134
rect 21062 614898 21146 615134
rect 21382 614898 21414 615134
rect 20794 579454 21414 614898
rect 20794 579218 20826 579454
rect 21062 579218 21146 579454
rect 21382 579218 21414 579454
rect 20794 579134 21414 579218
rect 20794 578898 20826 579134
rect 21062 578898 21146 579134
rect 21382 578898 21414 579134
rect 20794 543454 21414 578898
rect 20794 543218 20826 543454
rect 21062 543218 21146 543454
rect 21382 543218 21414 543454
rect 20794 543134 21414 543218
rect 20794 542898 20826 543134
rect 21062 542898 21146 543134
rect 21382 542898 21414 543134
rect 20794 507454 21414 542898
rect 20794 507218 20826 507454
rect 21062 507218 21146 507454
rect 21382 507218 21414 507454
rect 20794 507134 21414 507218
rect 20794 506898 20826 507134
rect 21062 506898 21146 507134
rect 21382 506898 21414 507134
rect 20794 471454 21414 506898
rect 20794 471218 20826 471454
rect 21062 471218 21146 471454
rect 21382 471218 21414 471454
rect 20794 471134 21414 471218
rect 20794 470898 20826 471134
rect 21062 470898 21146 471134
rect 21382 470898 21414 471134
rect 20794 435454 21414 470898
rect 20794 435218 20826 435454
rect 21062 435218 21146 435454
rect 21382 435218 21414 435454
rect 20794 435134 21414 435218
rect 20794 434898 20826 435134
rect 21062 434898 21146 435134
rect 21382 434898 21414 435134
rect 20794 399454 21414 434898
rect 20794 399218 20826 399454
rect 21062 399218 21146 399454
rect 21382 399218 21414 399454
rect 20794 399134 21414 399218
rect 20794 398898 20826 399134
rect 21062 398898 21146 399134
rect 21382 398898 21414 399134
rect 20794 363454 21414 398898
rect 20794 363218 20826 363454
rect 21062 363218 21146 363454
rect 21382 363218 21414 363454
rect 20794 363134 21414 363218
rect 20794 362898 20826 363134
rect 21062 362898 21146 363134
rect 21382 362898 21414 363134
rect 20794 327454 21414 362898
rect 20794 327218 20826 327454
rect 21062 327218 21146 327454
rect 21382 327218 21414 327454
rect 20794 327134 21414 327218
rect 20794 326898 20826 327134
rect 21062 326898 21146 327134
rect 21382 326898 21414 327134
rect 20794 291454 21414 326898
rect 20794 291218 20826 291454
rect 21062 291218 21146 291454
rect 21382 291218 21414 291454
rect 20794 291134 21414 291218
rect 20794 290898 20826 291134
rect 21062 290898 21146 291134
rect 21382 290898 21414 291134
rect 20794 255454 21414 290898
rect 20794 255218 20826 255454
rect 21062 255218 21146 255454
rect 21382 255218 21414 255454
rect 20794 255134 21414 255218
rect 20794 254898 20826 255134
rect 21062 254898 21146 255134
rect 21382 254898 21414 255134
rect 20794 219454 21414 254898
rect 20794 219218 20826 219454
rect 21062 219218 21146 219454
rect 21382 219218 21414 219454
rect 20794 219134 21414 219218
rect 20794 218898 20826 219134
rect 21062 218898 21146 219134
rect 21382 218898 21414 219134
rect 20794 183454 21414 218898
rect 20794 183218 20826 183454
rect 21062 183218 21146 183454
rect 21382 183218 21414 183454
rect 20794 183134 21414 183218
rect 20794 182898 20826 183134
rect 21062 182898 21146 183134
rect 21382 182898 21414 183134
rect 20794 147454 21414 182898
rect 20794 147218 20826 147454
rect 21062 147218 21146 147454
rect 21382 147218 21414 147454
rect 20794 147134 21414 147218
rect 20794 146898 20826 147134
rect 21062 146898 21146 147134
rect 21382 146898 21414 147134
rect 20794 111454 21414 146898
rect 20794 111218 20826 111454
rect 21062 111218 21146 111454
rect 21382 111218 21414 111454
rect 20794 111134 21414 111218
rect 20794 110898 20826 111134
rect 21062 110898 21146 111134
rect 21382 110898 21414 111134
rect 20794 75454 21414 110898
rect 20794 75218 20826 75454
rect 21062 75218 21146 75454
rect 21382 75218 21414 75454
rect 20794 75134 21414 75218
rect 20794 74898 20826 75134
rect 21062 74898 21146 75134
rect 21382 74898 21414 75134
rect 20794 74295 21414 74898
rect 21954 680614 22574 711002
rect 31954 710598 32574 711590
rect 31954 710362 31986 710598
rect 32222 710362 32306 710598
rect 32542 710362 32574 710598
rect 31954 710278 32574 710362
rect 31954 710042 31986 710278
rect 32222 710042 32306 710278
rect 32542 710042 32574 710278
rect 28234 708678 28854 709670
rect 28234 708442 28266 708678
rect 28502 708442 28586 708678
rect 28822 708442 28854 708678
rect 28234 708358 28854 708442
rect 28234 708122 28266 708358
rect 28502 708122 28586 708358
rect 28822 708122 28854 708358
rect 21954 680378 21986 680614
rect 22222 680378 22306 680614
rect 22542 680378 22574 680614
rect 21954 680294 22574 680378
rect 21954 680058 21986 680294
rect 22222 680058 22306 680294
rect 22542 680058 22574 680294
rect 21954 644614 22574 680058
rect 21954 644378 21986 644614
rect 22222 644378 22306 644614
rect 22542 644378 22574 644614
rect 21954 644294 22574 644378
rect 21954 644058 21986 644294
rect 22222 644058 22306 644294
rect 22542 644058 22574 644294
rect 21954 608614 22574 644058
rect 21954 608378 21986 608614
rect 22222 608378 22306 608614
rect 22542 608378 22574 608614
rect 21954 608294 22574 608378
rect 21954 608058 21986 608294
rect 22222 608058 22306 608294
rect 22542 608058 22574 608294
rect 21954 572614 22574 608058
rect 21954 572378 21986 572614
rect 22222 572378 22306 572614
rect 22542 572378 22574 572614
rect 21954 572294 22574 572378
rect 21954 572058 21986 572294
rect 22222 572058 22306 572294
rect 22542 572058 22574 572294
rect 21954 536614 22574 572058
rect 21954 536378 21986 536614
rect 22222 536378 22306 536614
rect 22542 536378 22574 536614
rect 21954 536294 22574 536378
rect 21954 536058 21986 536294
rect 22222 536058 22306 536294
rect 22542 536058 22574 536294
rect 21954 500614 22574 536058
rect 21954 500378 21986 500614
rect 22222 500378 22306 500614
rect 22542 500378 22574 500614
rect 21954 500294 22574 500378
rect 21954 500058 21986 500294
rect 22222 500058 22306 500294
rect 22542 500058 22574 500294
rect 21954 464614 22574 500058
rect 21954 464378 21986 464614
rect 22222 464378 22306 464614
rect 22542 464378 22574 464614
rect 21954 464294 22574 464378
rect 21954 464058 21986 464294
rect 22222 464058 22306 464294
rect 22542 464058 22574 464294
rect 21954 428614 22574 464058
rect 21954 428378 21986 428614
rect 22222 428378 22306 428614
rect 22542 428378 22574 428614
rect 21954 428294 22574 428378
rect 21954 428058 21986 428294
rect 22222 428058 22306 428294
rect 22542 428058 22574 428294
rect 21954 392614 22574 428058
rect 21954 392378 21986 392614
rect 22222 392378 22306 392614
rect 22542 392378 22574 392614
rect 21954 392294 22574 392378
rect 21954 392058 21986 392294
rect 22222 392058 22306 392294
rect 22542 392058 22574 392294
rect 21954 356614 22574 392058
rect 21954 356378 21986 356614
rect 22222 356378 22306 356614
rect 22542 356378 22574 356614
rect 21954 356294 22574 356378
rect 21954 356058 21986 356294
rect 22222 356058 22306 356294
rect 22542 356058 22574 356294
rect 21954 320614 22574 356058
rect 21954 320378 21986 320614
rect 22222 320378 22306 320614
rect 22542 320378 22574 320614
rect 21954 320294 22574 320378
rect 21954 320058 21986 320294
rect 22222 320058 22306 320294
rect 22542 320058 22574 320294
rect 21954 284614 22574 320058
rect 21954 284378 21986 284614
rect 22222 284378 22306 284614
rect 22542 284378 22574 284614
rect 21954 284294 22574 284378
rect 21954 284058 21986 284294
rect 22222 284058 22306 284294
rect 22542 284058 22574 284294
rect 21954 248614 22574 284058
rect 21954 248378 21986 248614
rect 22222 248378 22306 248614
rect 22542 248378 22574 248614
rect 21954 248294 22574 248378
rect 21954 248058 21986 248294
rect 22222 248058 22306 248294
rect 22542 248058 22574 248294
rect 21954 212614 22574 248058
rect 21954 212378 21986 212614
rect 22222 212378 22306 212614
rect 22542 212378 22574 212614
rect 21954 212294 22574 212378
rect 21954 212058 21986 212294
rect 22222 212058 22306 212294
rect 22542 212058 22574 212294
rect 21954 176614 22574 212058
rect 21954 176378 21986 176614
rect 22222 176378 22306 176614
rect 22542 176378 22574 176614
rect 21954 176294 22574 176378
rect 21954 176058 21986 176294
rect 22222 176058 22306 176294
rect 22542 176058 22574 176294
rect 21954 140614 22574 176058
rect 21954 140378 21986 140614
rect 22222 140378 22306 140614
rect 22542 140378 22574 140614
rect 21954 140294 22574 140378
rect 21954 140058 21986 140294
rect 22222 140058 22306 140294
rect 22542 140058 22574 140294
rect 21954 104614 22574 140058
rect 21954 104378 21986 104614
rect 22222 104378 22306 104614
rect 22542 104378 22574 104614
rect 21954 104294 22574 104378
rect 21954 104058 21986 104294
rect 22222 104058 22306 104294
rect 22542 104058 22574 104294
rect 21954 74295 22574 104058
rect 24514 706758 25134 707750
rect 24514 706522 24546 706758
rect 24782 706522 24866 706758
rect 25102 706522 25134 706758
rect 24514 706438 25134 706522
rect 24514 706202 24546 706438
rect 24782 706202 24866 706438
rect 25102 706202 25134 706438
rect 24514 691174 25134 706202
rect 24514 690938 24546 691174
rect 24782 690938 24866 691174
rect 25102 690938 25134 691174
rect 24514 690854 25134 690938
rect 24514 690618 24546 690854
rect 24782 690618 24866 690854
rect 25102 690618 25134 690854
rect 24514 655174 25134 690618
rect 24514 654938 24546 655174
rect 24782 654938 24866 655174
rect 25102 654938 25134 655174
rect 24514 654854 25134 654938
rect 24514 654618 24546 654854
rect 24782 654618 24866 654854
rect 25102 654618 25134 654854
rect 24514 619174 25134 654618
rect 24514 618938 24546 619174
rect 24782 618938 24866 619174
rect 25102 618938 25134 619174
rect 24514 618854 25134 618938
rect 24514 618618 24546 618854
rect 24782 618618 24866 618854
rect 25102 618618 25134 618854
rect 24514 583174 25134 618618
rect 24514 582938 24546 583174
rect 24782 582938 24866 583174
rect 25102 582938 25134 583174
rect 24514 582854 25134 582938
rect 24514 582618 24546 582854
rect 24782 582618 24866 582854
rect 25102 582618 25134 582854
rect 24514 547174 25134 582618
rect 24514 546938 24546 547174
rect 24782 546938 24866 547174
rect 25102 546938 25134 547174
rect 24514 546854 25134 546938
rect 24514 546618 24546 546854
rect 24782 546618 24866 546854
rect 25102 546618 25134 546854
rect 24514 511174 25134 546618
rect 24514 510938 24546 511174
rect 24782 510938 24866 511174
rect 25102 510938 25134 511174
rect 24514 510854 25134 510938
rect 24514 510618 24546 510854
rect 24782 510618 24866 510854
rect 25102 510618 25134 510854
rect 24514 475174 25134 510618
rect 24514 474938 24546 475174
rect 24782 474938 24866 475174
rect 25102 474938 25134 475174
rect 24514 474854 25134 474938
rect 24514 474618 24546 474854
rect 24782 474618 24866 474854
rect 25102 474618 25134 474854
rect 24514 439174 25134 474618
rect 24514 438938 24546 439174
rect 24782 438938 24866 439174
rect 25102 438938 25134 439174
rect 24514 438854 25134 438938
rect 24514 438618 24546 438854
rect 24782 438618 24866 438854
rect 25102 438618 25134 438854
rect 24514 403174 25134 438618
rect 24514 402938 24546 403174
rect 24782 402938 24866 403174
rect 25102 402938 25134 403174
rect 24514 402854 25134 402938
rect 24514 402618 24546 402854
rect 24782 402618 24866 402854
rect 25102 402618 25134 402854
rect 24514 367174 25134 402618
rect 24514 366938 24546 367174
rect 24782 366938 24866 367174
rect 25102 366938 25134 367174
rect 24514 366854 25134 366938
rect 24514 366618 24546 366854
rect 24782 366618 24866 366854
rect 25102 366618 25134 366854
rect 24514 331174 25134 366618
rect 24514 330938 24546 331174
rect 24782 330938 24866 331174
rect 25102 330938 25134 331174
rect 24514 330854 25134 330938
rect 24514 330618 24546 330854
rect 24782 330618 24866 330854
rect 25102 330618 25134 330854
rect 24514 295174 25134 330618
rect 24514 294938 24546 295174
rect 24782 294938 24866 295174
rect 25102 294938 25134 295174
rect 24514 294854 25134 294938
rect 24514 294618 24546 294854
rect 24782 294618 24866 294854
rect 25102 294618 25134 294854
rect 24514 259174 25134 294618
rect 24514 258938 24546 259174
rect 24782 258938 24866 259174
rect 25102 258938 25134 259174
rect 24514 258854 25134 258938
rect 24514 258618 24546 258854
rect 24782 258618 24866 258854
rect 25102 258618 25134 258854
rect 24514 223174 25134 258618
rect 24514 222938 24546 223174
rect 24782 222938 24866 223174
rect 25102 222938 25134 223174
rect 24514 222854 25134 222938
rect 24514 222618 24546 222854
rect 24782 222618 24866 222854
rect 25102 222618 25134 222854
rect 24514 187174 25134 222618
rect 24514 186938 24546 187174
rect 24782 186938 24866 187174
rect 25102 186938 25134 187174
rect 24514 186854 25134 186938
rect 24514 186618 24546 186854
rect 24782 186618 24866 186854
rect 25102 186618 25134 186854
rect 24514 151174 25134 186618
rect 24514 150938 24546 151174
rect 24782 150938 24866 151174
rect 25102 150938 25134 151174
rect 24514 150854 25134 150938
rect 24514 150618 24546 150854
rect 24782 150618 24866 150854
rect 25102 150618 25134 150854
rect 24514 115174 25134 150618
rect 24514 114938 24546 115174
rect 24782 114938 24866 115174
rect 25102 114938 25134 115174
rect 24514 114854 25134 114938
rect 24514 114618 24546 114854
rect 24782 114618 24866 114854
rect 25102 114618 25134 114854
rect 24514 79174 25134 114618
rect 24514 78938 24546 79174
rect 24782 78938 24866 79174
rect 25102 78938 25134 79174
rect 24514 78854 25134 78938
rect 24514 78618 24546 78854
rect 24782 78618 24866 78854
rect 25102 78618 25134 78854
rect 24514 74295 25134 78618
rect 28234 694894 28854 708122
rect 28234 694658 28266 694894
rect 28502 694658 28586 694894
rect 28822 694658 28854 694894
rect 28234 694574 28854 694658
rect 28234 694338 28266 694574
rect 28502 694338 28586 694574
rect 28822 694338 28854 694574
rect 28234 658894 28854 694338
rect 28234 658658 28266 658894
rect 28502 658658 28586 658894
rect 28822 658658 28854 658894
rect 28234 658574 28854 658658
rect 28234 658338 28266 658574
rect 28502 658338 28586 658574
rect 28822 658338 28854 658574
rect 28234 622894 28854 658338
rect 28234 622658 28266 622894
rect 28502 622658 28586 622894
rect 28822 622658 28854 622894
rect 28234 622574 28854 622658
rect 28234 622338 28266 622574
rect 28502 622338 28586 622574
rect 28822 622338 28854 622574
rect 28234 586894 28854 622338
rect 28234 586658 28266 586894
rect 28502 586658 28586 586894
rect 28822 586658 28854 586894
rect 28234 586574 28854 586658
rect 28234 586338 28266 586574
rect 28502 586338 28586 586574
rect 28822 586338 28854 586574
rect 28234 550894 28854 586338
rect 28234 550658 28266 550894
rect 28502 550658 28586 550894
rect 28822 550658 28854 550894
rect 28234 550574 28854 550658
rect 28234 550338 28266 550574
rect 28502 550338 28586 550574
rect 28822 550338 28854 550574
rect 28234 514894 28854 550338
rect 28234 514658 28266 514894
rect 28502 514658 28586 514894
rect 28822 514658 28854 514894
rect 28234 514574 28854 514658
rect 28234 514338 28266 514574
rect 28502 514338 28586 514574
rect 28822 514338 28854 514574
rect 28234 478894 28854 514338
rect 28234 478658 28266 478894
rect 28502 478658 28586 478894
rect 28822 478658 28854 478894
rect 28234 478574 28854 478658
rect 28234 478338 28266 478574
rect 28502 478338 28586 478574
rect 28822 478338 28854 478574
rect 28234 442894 28854 478338
rect 28234 442658 28266 442894
rect 28502 442658 28586 442894
rect 28822 442658 28854 442894
rect 28234 442574 28854 442658
rect 28234 442338 28266 442574
rect 28502 442338 28586 442574
rect 28822 442338 28854 442574
rect 28234 406894 28854 442338
rect 28234 406658 28266 406894
rect 28502 406658 28586 406894
rect 28822 406658 28854 406894
rect 28234 406574 28854 406658
rect 28234 406338 28266 406574
rect 28502 406338 28586 406574
rect 28822 406338 28854 406574
rect 28234 370894 28854 406338
rect 28234 370658 28266 370894
rect 28502 370658 28586 370894
rect 28822 370658 28854 370894
rect 28234 370574 28854 370658
rect 28234 370338 28266 370574
rect 28502 370338 28586 370574
rect 28822 370338 28854 370574
rect 28234 334894 28854 370338
rect 28234 334658 28266 334894
rect 28502 334658 28586 334894
rect 28822 334658 28854 334894
rect 28234 334574 28854 334658
rect 28234 334338 28266 334574
rect 28502 334338 28586 334574
rect 28822 334338 28854 334574
rect 28234 298894 28854 334338
rect 28234 298658 28266 298894
rect 28502 298658 28586 298894
rect 28822 298658 28854 298894
rect 28234 298574 28854 298658
rect 28234 298338 28266 298574
rect 28502 298338 28586 298574
rect 28822 298338 28854 298574
rect 28234 262894 28854 298338
rect 28234 262658 28266 262894
rect 28502 262658 28586 262894
rect 28822 262658 28854 262894
rect 28234 262574 28854 262658
rect 28234 262338 28266 262574
rect 28502 262338 28586 262574
rect 28822 262338 28854 262574
rect 28234 226894 28854 262338
rect 28234 226658 28266 226894
rect 28502 226658 28586 226894
rect 28822 226658 28854 226894
rect 28234 226574 28854 226658
rect 28234 226338 28266 226574
rect 28502 226338 28586 226574
rect 28822 226338 28854 226574
rect 28234 190894 28854 226338
rect 28234 190658 28266 190894
rect 28502 190658 28586 190894
rect 28822 190658 28854 190894
rect 28234 190574 28854 190658
rect 28234 190338 28266 190574
rect 28502 190338 28586 190574
rect 28822 190338 28854 190574
rect 28234 154894 28854 190338
rect 28234 154658 28266 154894
rect 28502 154658 28586 154894
rect 28822 154658 28854 154894
rect 28234 154574 28854 154658
rect 28234 154338 28266 154574
rect 28502 154338 28586 154574
rect 28822 154338 28854 154574
rect 28234 118894 28854 154338
rect 28234 118658 28266 118894
rect 28502 118658 28586 118894
rect 28822 118658 28854 118894
rect 28234 118574 28854 118658
rect 28234 118338 28266 118574
rect 28502 118338 28586 118574
rect 28822 118338 28854 118574
rect 28234 82894 28854 118338
rect 28234 82658 28266 82894
rect 28502 82658 28586 82894
rect 28822 82658 28854 82894
rect 28234 82574 28854 82658
rect 28234 82338 28266 82574
rect 28502 82338 28586 82574
rect 28822 82338 28854 82574
rect 28234 74295 28854 82338
rect 30794 705798 31414 705830
rect 30794 705562 30826 705798
rect 31062 705562 31146 705798
rect 31382 705562 31414 705798
rect 30794 705478 31414 705562
rect 30794 705242 30826 705478
rect 31062 705242 31146 705478
rect 31382 705242 31414 705478
rect 30794 669454 31414 705242
rect 30794 669218 30826 669454
rect 31062 669218 31146 669454
rect 31382 669218 31414 669454
rect 30794 669134 31414 669218
rect 30794 668898 30826 669134
rect 31062 668898 31146 669134
rect 31382 668898 31414 669134
rect 30794 633454 31414 668898
rect 30794 633218 30826 633454
rect 31062 633218 31146 633454
rect 31382 633218 31414 633454
rect 30794 633134 31414 633218
rect 30794 632898 30826 633134
rect 31062 632898 31146 633134
rect 31382 632898 31414 633134
rect 30794 597454 31414 632898
rect 30794 597218 30826 597454
rect 31062 597218 31146 597454
rect 31382 597218 31414 597454
rect 30794 597134 31414 597218
rect 30794 596898 30826 597134
rect 31062 596898 31146 597134
rect 31382 596898 31414 597134
rect 30794 561454 31414 596898
rect 30794 561218 30826 561454
rect 31062 561218 31146 561454
rect 31382 561218 31414 561454
rect 30794 561134 31414 561218
rect 30794 560898 30826 561134
rect 31062 560898 31146 561134
rect 31382 560898 31414 561134
rect 30794 525454 31414 560898
rect 30794 525218 30826 525454
rect 31062 525218 31146 525454
rect 31382 525218 31414 525454
rect 30794 525134 31414 525218
rect 30794 524898 30826 525134
rect 31062 524898 31146 525134
rect 31382 524898 31414 525134
rect 30794 489454 31414 524898
rect 30794 489218 30826 489454
rect 31062 489218 31146 489454
rect 31382 489218 31414 489454
rect 30794 489134 31414 489218
rect 30794 488898 30826 489134
rect 31062 488898 31146 489134
rect 31382 488898 31414 489134
rect 30794 453454 31414 488898
rect 30794 453218 30826 453454
rect 31062 453218 31146 453454
rect 31382 453218 31414 453454
rect 30794 453134 31414 453218
rect 30794 452898 30826 453134
rect 31062 452898 31146 453134
rect 31382 452898 31414 453134
rect 30794 417454 31414 452898
rect 30794 417218 30826 417454
rect 31062 417218 31146 417454
rect 31382 417218 31414 417454
rect 30794 417134 31414 417218
rect 30794 416898 30826 417134
rect 31062 416898 31146 417134
rect 31382 416898 31414 417134
rect 30794 381454 31414 416898
rect 30794 381218 30826 381454
rect 31062 381218 31146 381454
rect 31382 381218 31414 381454
rect 30794 381134 31414 381218
rect 30794 380898 30826 381134
rect 31062 380898 31146 381134
rect 31382 380898 31414 381134
rect 30794 345454 31414 380898
rect 30794 345218 30826 345454
rect 31062 345218 31146 345454
rect 31382 345218 31414 345454
rect 30794 345134 31414 345218
rect 30794 344898 30826 345134
rect 31062 344898 31146 345134
rect 31382 344898 31414 345134
rect 30794 309454 31414 344898
rect 30794 309218 30826 309454
rect 31062 309218 31146 309454
rect 31382 309218 31414 309454
rect 30794 309134 31414 309218
rect 30794 308898 30826 309134
rect 31062 308898 31146 309134
rect 31382 308898 31414 309134
rect 30794 273454 31414 308898
rect 30794 273218 30826 273454
rect 31062 273218 31146 273454
rect 31382 273218 31414 273454
rect 30794 273134 31414 273218
rect 30794 272898 30826 273134
rect 31062 272898 31146 273134
rect 31382 272898 31414 273134
rect 30794 237454 31414 272898
rect 30794 237218 30826 237454
rect 31062 237218 31146 237454
rect 31382 237218 31414 237454
rect 30794 237134 31414 237218
rect 30794 236898 30826 237134
rect 31062 236898 31146 237134
rect 31382 236898 31414 237134
rect 30794 201454 31414 236898
rect 30794 201218 30826 201454
rect 31062 201218 31146 201454
rect 31382 201218 31414 201454
rect 30794 201134 31414 201218
rect 30794 200898 30826 201134
rect 31062 200898 31146 201134
rect 31382 200898 31414 201134
rect 30794 165454 31414 200898
rect 30794 165218 30826 165454
rect 31062 165218 31146 165454
rect 31382 165218 31414 165454
rect 30794 165134 31414 165218
rect 30794 164898 30826 165134
rect 31062 164898 31146 165134
rect 31382 164898 31414 165134
rect 30794 129454 31414 164898
rect 30794 129218 30826 129454
rect 31062 129218 31146 129454
rect 31382 129218 31414 129454
rect 30794 129134 31414 129218
rect 30794 128898 30826 129134
rect 31062 128898 31146 129134
rect 31382 128898 31414 129134
rect 30794 93454 31414 128898
rect 30794 93218 30826 93454
rect 31062 93218 31146 93454
rect 31382 93218 31414 93454
rect 30794 93134 31414 93218
rect 30794 92898 30826 93134
rect 31062 92898 31146 93134
rect 31382 92898 31414 93134
rect 30794 74295 31414 92898
rect 31954 698614 32574 710042
rect 41954 711558 42574 711590
rect 41954 711322 41986 711558
rect 42222 711322 42306 711558
rect 42542 711322 42574 711558
rect 41954 711238 42574 711322
rect 41954 711002 41986 711238
rect 42222 711002 42306 711238
rect 42542 711002 42574 711238
rect 38234 709638 38854 709670
rect 38234 709402 38266 709638
rect 38502 709402 38586 709638
rect 38822 709402 38854 709638
rect 38234 709318 38854 709402
rect 38234 709082 38266 709318
rect 38502 709082 38586 709318
rect 38822 709082 38854 709318
rect 31954 698378 31986 698614
rect 32222 698378 32306 698614
rect 32542 698378 32574 698614
rect 31954 698294 32574 698378
rect 31954 698058 31986 698294
rect 32222 698058 32306 698294
rect 32542 698058 32574 698294
rect 31954 662614 32574 698058
rect 31954 662378 31986 662614
rect 32222 662378 32306 662614
rect 32542 662378 32574 662614
rect 31954 662294 32574 662378
rect 31954 662058 31986 662294
rect 32222 662058 32306 662294
rect 32542 662058 32574 662294
rect 31954 626614 32574 662058
rect 31954 626378 31986 626614
rect 32222 626378 32306 626614
rect 32542 626378 32574 626614
rect 31954 626294 32574 626378
rect 31954 626058 31986 626294
rect 32222 626058 32306 626294
rect 32542 626058 32574 626294
rect 31954 590614 32574 626058
rect 31954 590378 31986 590614
rect 32222 590378 32306 590614
rect 32542 590378 32574 590614
rect 31954 590294 32574 590378
rect 31954 590058 31986 590294
rect 32222 590058 32306 590294
rect 32542 590058 32574 590294
rect 31954 554614 32574 590058
rect 31954 554378 31986 554614
rect 32222 554378 32306 554614
rect 32542 554378 32574 554614
rect 31954 554294 32574 554378
rect 31954 554058 31986 554294
rect 32222 554058 32306 554294
rect 32542 554058 32574 554294
rect 31954 518614 32574 554058
rect 31954 518378 31986 518614
rect 32222 518378 32306 518614
rect 32542 518378 32574 518614
rect 31954 518294 32574 518378
rect 31954 518058 31986 518294
rect 32222 518058 32306 518294
rect 32542 518058 32574 518294
rect 31954 482614 32574 518058
rect 31954 482378 31986 482614
rect 32222 482378 32306 482614
rect 32542 482378 32574 482614
rect 31954 482294 32574 482378
rect 31954 482058 31986 482294
rect 32222 482058 32306 482294
rect 32542 482058 32574 482294
rect 31954 446614 32574 482058
rect 31954 446378 31986 446614
rect 32222 446378 32306 446614
rect 32542 446378 32574 446614
rect 31954 446294 32574 446378
rect 31954 446058 31986 446294
rect 32222 446058 32306 446294
rect 32542 446058 32574 446294
rect 31954 410614 32574 446058
rect 31954 410378 31986 410614
rect 32222 410378 32306 410614
rect 32542 410378 32574 410614
rect 31954 410294 32574 410378
rect 31954 410058 31986 410294
rect 32222 410058 32306 410294
rect 32542 410058 32574 410294
rect 31954 374614 32574 410058
rect 31954 374378 31986 374614
rect 32222 374378 32306 374614
rect 32542 374378 32574 374614
rect 31954 374294 32574 374378
rect 31954 374058 31986 374294
rect 32222 374058 32306 374294
rect 32542 374058 32574 374294
rect 31954 338614 32574 374058
rect 31954 338378 31986 338614
rect 32222 338378 32306 338614
rect 32542 338378 32574 338614
rect 31954 338294 32574 338378
rect 31954 338058 31986 338294
rect 32222 338058 32306 338294
rect 32542 338058 32574 338294
rect 31954 302614 32574 338058
rect 31954 302378 31986 302614
rect 32222 302378 32306 302614
rect 32542 302378 32574 302614
rect 31954 302294 32574 302378
rect 31954 302058 31986 302294
rect 32222 302058 32306 302294
rect 32542 302058 32574 302294
rect 31954 266614 32574 302058
rect 31954 266378 31986 266614
rect 32222 266378 32306 266614
rect 32542 266378 32574 266614
rect 31954 266294 32574 266378
rect 31954 266058 31986 266294
rect 32222 266058 32306 266294
rect 32542 266058 32574 266294
rect 31954 230614 32574 266058
rect 31954 230378 31986 230614
rect 32222 230378 32306 230614
rect 32542 230378 32574 230614
rect 31954 230294 32574 230378
rect 31954 230058 31986 230294
rect 32222 230058 32306 230294
rect 32542 230058 32574 230294
rect 31954 194614 32574 230058
rect 31954 194378 31986 194614
rect 32222 194378 32306 194614
rect 32542 194378 32574 194614
rect 31954 194294 32574 194378
rect 31954 194058 31986 194294
rect 32222 194058 32306 194294
rect 32542 194058 32574 194294
rect 31954 158614 32574 194058
rect 31954 158378 31986 158614
rect 32222 158378 32306 158614
rect 32542 158378 32574 158614
rect 31954 158294 32574 158378
rect 31954 158058 31986 158294
rect 32222 158058 32306 158294
rect 32542 158058 32574 158294
rect 31954 122614 32574 158058
rect 31954 122378 31986 122614
rect 32222 122378 32306 122614
rect 32542 122378 32574 122614
rect 31954 122294 32574 122378
rect 31954 122058 31986 122294
rect 32222 122058 32306 122294
rect 32542 122058 32574 122294
rect 31954 86614 32574 122058
rect 31954 86378 31986 86614
rect 32222 86378 32306 86614
rect 32542 86378 32574 86614
rect 31954 86294 32574 86378
rect 31954 86058 31986 86294
rect 32222 86058 32306 86294
rect 32542 86058 32574 86294
rect 31954 74295 32574 86058
rect 34514 707718 35134 707750
rect 34514 707482 34546 707718
rect 34782 707482 34866 707718
rect 35102 707482 35134 707718
rect 34514 707398 35134 707482
rect 34514 707162 34546 707398
rect 34782 707162 34866 707398
rect 35102 707162 35134 707398
rect 34514 673174 35134 707162
rect 34514 672938 34546 673174
rect 34782 672938 34866 673174
rect 35102 672938 35134 673174
rect 34514 672854 35134 672938
rect 34514 672618 34546 672854
rect 34782 672618 34866 672854
rect 35102 672618 35134 672854
rect 34514 637174 35134 672618
rect 34514 636938 34546 637174
rect 34782 636938 34866 637174
rect 35102 636938 35134 637174
rect 34514 636854 35134 636938
rect 34514 636618 34546 636854
rect 34782 636618 34866 636854
rect 35102 636618 35134 636854
rect 34514 601174 35134 636618
rect 34514 600938 34546 601174
rect 34782 600938 34866 601174
rect 35102 600938 35134 601174
rect 34514 600854 35134 600938
rect 34514 600618 34546 600854
rect 34782 600618 34866 600854
rect 35102 600618 35134 600854
rect 34514 565174 35134 600618
rect 34514 564938 34546 565174
rect 34782 564938 34866 565174
rect 35102 564938 35134 565174
rect 34514 564854 35134 564938
rect 34514 564618 34546 564854
rect 34782 564618 34866 564854
rect 35102 564618 35134 564854
rect 34514 529174 35134 564618
rect 34514 528938 34546 529174
rect 34782 528938 34866 529174
rect 35102 528938 35134 529174
rect 34514 528854 35134 528938
rect 34514 528618 34546 528854
rect 34782 528618 34866 528854
rect 35102 528618 35134 528854
rect 34514 493174 35134 528618
rect 34514 492938 34546 493174
rect 34782 492938 34866 493174
rect 35102 492938 35134 493174
rect 34514 492854 35134 492938
rect 34514 492618 34546 492854
rect 34782 492618 34866 492854
rect 35102 492618 35134 492854
rect 34514 457174 35134 492618
rect 34514 456938 34546 457174
rect 34782 456938 34866 457174
rect 35102 456938 35134 457174
rect 34514 456854 35134 456938
rect 34514 456618 34546 456854
rect 34782 456618 34866 456854
rect 35102 456618 35134 456854
rect 34514 421174 35134 456618
rect 34514 420938 34546 421174
rect 34782 420938 34866 421174
rect 35102 420938 35134 421174
rect 34514 420854 35134 420938
rect 34514 420618 34546 420854
rect 34782 420618 34866 420854
rect 35102 420618 35134 420854
rect 34514 385174 35134 420618
rect 34514 384938 34546 385174
rect 34782 384938 34866 385174
rect 35102 384938 35134 385174
rect 34514 384854 35134 384938
rect 34514 384618 34546 384854
rect 34782 384618 34866 384854
rect 35102 384618 35134 384854
rect 34514 349174 35134 384618
rect 34514 348938 34546 349174
rect 34782 348938 34866 349174
rect 35102 348938 35134 349174
rect 34514 348854 35134 348938
rect 34514 348618 34546 348854
rect 34782 348618 34866 348854
rect 35102 348618 35134 348854
rect 34514 313174 35134 348618
rect 34514 312938 34546 313174
rect 34782 312938 34866 313174
rect 35102 312938 35134 313174
rect 34514 312854 35134 312938
rect 34514 312618 34546 312854
rect 34782 312618 34866 312854
rect 35102 312618 35134 312854
rect 34514 277174 35134 312618
rect 34514 276938 34546 277174
rect 34782 276938 34866 277174
rect 35102 276938 35134 277174
rect 34514 276854 35134 276938
rect 34514 276618 34546 276854
rect 34782 276618 34866 276854
rect 35102 276618 35134 276854
rect 34514 241174 35134 276618
rect 34514 240938 34546 241174
rect 34782 240938 34866 241174
rect 35102 240938 35134 241174
rect 34514 240854 35134 240938
rect 34514 240618 34546 240854
rect 34782 240618 34866 240854
rect 35102 240618 35134 240854
rect 34514 205174 35134 240618
rect 34514 204938 34546 205174
rect 34782 204938 34866 205174
rect 35102 204938 35134 205174
rect 34514 204854 35134 204938
rect 34514 204618 34546 204854
rect 34782 204618 34866 204854
rect 35102 204618 35134 204854
rect 34514 169174 35134 204618
rect 34514 168938 34546 169174
rect 34782 168938 34866 169174
rect 35102 168938 35134 169174
rect 34514 168854 35134 168938
rect 34514 168618 34546 168854
rect 34782 168618 34866 168854
rect 35102 168618 35134 168854
rect 34514 133174 35134 168618
rect 34514 132938 34546 133174
rect 34782 132938 34866 133174
rect 35102 132938 35134 133174
rect 34514 132854 35134 132938
rect 34514 132618 34546 132854
rect 34782 132618 34866 132854
rect 35102 132618 35134 132854
rect 34514 97174 35134 132618
rect 34514 96938 34546 97174
rect 34782 96938 34866 97174
rect 35102 96938 35134 97174
rect 34514 96854 35134 96938
rect 34514 96618 34546 96854
rect 34782 96618 34866 96854
rect 35102 96618 35134 96854
rect 34514 74295 35134 96618
rect 38234 676894 38854 709082
rect 38234 676658 38266 676894
rect 38502 676658 38586 676894
rect 38822 676658 38854 676894
rect 38234 676574 38854 676658
rect 38234 676338 38266 676574
rect 38502 676338 38586 676574
rect 38822 676338 38854 676574
rect 38234 640894 38854 676338
rect 38234 640658 38266 640894
rect 38502 640658 38586 640894
rect 38822 640658 38854 640894
rect 38234 640574 38854 640658
rect 38234 640338 38266 640574
rect 38502 640338 38586 640574
rect 38822 640338 38854 640574
rect 38234 604894 38854 640338
rect 38234 604658 38266 604894
rect 38502 604658 38586 604894
rect 38822 604658 38854 604894
rect 38234 604574 38854 604658
rect 38234 604338 38266 604574
rect 38502 604338 38586 604574
rect 38822 604338 38854 604574
rect 38234 568894 38854 604338
rect 38234 568658 38266 568894
rect 38502 568658 38586 568894
rect 38822 568658 38854 568894
rect 38234 568574 38854 568658
rect 38234 568338 38266 568574
rect 38502 568338 38586 568574
rect 38822 568338 38854 568574
rect 38234 532894 38854 568338
rect 38234 532658 38266 532894
rect 38502 532658 38586 532894
rect 38822 532658 38854 532894
rect 38234 532574 38854 532658
rect 38234 532338 38266 532574
rect 38502 532338 38586 532574
rect 38822 532338 38854 532574
rect 38234 496894 38854 532338
rect 38234 496658 38266 496894
rect 38502 496658 38586 496894
rect 38822 496658 38854 496894
rect 38234 496574 38854 496658
rect 38234 496338 38266 496574
rect 38502 496338 38586 496574
rect 38822 496338 38854 496574
rect 38234 460894 38854 496338
rect 38234 460658 38266 460894
rect 38502 460658 38586 460894
rect 38822 460658 38854 460894
rect 38234 460574 38854 460658
rect 38234 460338 38266 460574
rect 38502 460338 38586 460574
rect 38822 460338 38854 460574
rect 38234 424894 38854 460338
rect 38234 424658 38266 424894
rect 38502 424658 38586 424894
rect 38822 424658 38854 424894
rect 38234 424574 38854 424658
rect 38234 424338 38266 424574
rect 38502 424338 38586 424574
rect 38822 424338 38854 424574
rect 38234 388894 38854 424338
rect 38234 388658 38266 388894
rect 38502 388658 38586 388894
rect 38822 388658 38854 388894
rect 38234 388574 38854 388658
rect 38234 388338 38266 388574
rect 38502 388338 38586 388574
rect 38822 388338 38854 388574
rect 38234 352894 38854 388338
rect 38234 352658 38266 352894
rect 38502 352658 38586 352894
rect 38822 352658 38854 352894
rect 38234 352574 38854 352658
rect 38234 352338 38266 352574
rect 38502 352338 38586 352574
rect 38822 352338 38854 352574
rect 38234 316894 38854 352338
rect 38234 316658 38266 316894
rect 38502 316658 38586 316894
rect 38822 316658 38854 316894
rect 38234 316574 38854 316658
rect 38234 316338 38266 316574
rect 38502 316338 38586 316574
rect 38822 316338 38854 316574
rect 38234 280894 38854 316338
rect 38234 280658 38266 280894
rect 38502 280658 38586 280894
rect 38822 280658 38854 280894
rect 38234 280574 38854 280658
rect 38234 280338 38266 280574
rect 38502 280338 38586 280574
rect 38822 280338 38854 280574
rect 38234 244894 38854 280338
rect 38234 244658 38266 244894
rect 38502 244658 38586 244894
rect 38822 244658 38854 244894
rect 38234 244574 38854 244658
rect 38234 244338 38266 244574
rect 38502 244338 38586 244574
rect 38822 244338 38854 244574
rect 38234 208894 38854 244338
rect 38234 208658 38266 208894
rect 38502 208658 38586 208894
rect 38822 208658 38854 208894
rect 38234 208574 38854 208658
rect 38234 208338 38266 208574
rect 38502 208338 38586 208574
rect 38822 208338 38854 208574
rect 38234 172894 38854 208338
rect 38234 172658 38266 172894
rect 38502 172658 38586 172894
rect 38822 172658 38854 172894
rect 38234 172574 38854 172658
rect 38234 172338 38266 172574
rect 38502 172338 38586 172574
rect 38822 172338 38854 172574
rect 38234 136894 38854 172338
rect 38234 136658 38266 136894
rect 38502 136658 38586 136894
rect 38822 136658 38854 136894
rect 38234 136574 38854 136658
rect 38234 136338 38266 136574
rect 38502 136338 38586 136574
rect 38822 136338 38854 136574
rect 38234 100894 38854 136338
rect 38234 100658 38266 100894
rect 38502 100658 38586 100894
rect 38822 100658 38854 100894
rect 38234 100574 38854 100658
rect 38234 100338 38266 100574
rect 38502 100338 38586 100574
rect 38822 100338 38854 100574
rect 38234 74295 38854 100338
rect 40794 704838 41414 705830
rect 40794 704602 40826 704838
rect 41062 704602 41146 704838
rect 41382 704602 41414 704838
rect 40794 704518 41414 704602
rect 40794 704282 40826 704518
rect 41062 704282 41146 704518
rect 41382 704282 41414 704518
rect 40794 687454 41414 704282
rect 40794 687218 40826 687454
rect 41062 687218 41146 687454
rect 41382 687218 41414 687454
rect 40794 687134 41414 687218
rect 40794 686898 40826 687134
rect 41062 686898 41146 687134
rect 41382 686898 41414 687134
rect 40794 651454 41414 686898
rect 40794 651218 40826 651454
rect 41062 651218 41146 651454
rect 41382 651218 41414 651454
rect 40794 651134 41414 651218
rect 40794 650898 40826 651134
rect 41062 650898 41146 651134
rect 41382 650898 41414 651134
rect 40794 615454 41414 650898
rect 40794 615218 40826 615454
rect 41062 615218 41146 615454
rect 41382 615218 41414 615454
rect 40794 615134 41414 615218
rect 40794 614898 40826 615134
rect 41062 614898 41146 615134
rect 41382 614898 41414 615134
rect 40794 579454 41414 614898
rect 40794 579218 40826 579454
rect 41062 579218 41146 579454
rect 41382 579218 41414 579454
rect 40794 579134 41414 579218
rect 40794 578898 40826 579134
rect 41062 578898 41146 579134
rect 41382 578898 41414 579134
rect 40794 543454 41414 578898
rect 40794 543218 40826 543454
rect 41062 543218 41146 543454
rect 41382 543218 41414 543454
rect 40794 543134 41414 543218
rect 40794 542898 40826 543134
rect 41062 542898 41146 543134
rect 41382 542898 41414 543134
rect 40794 507454 41414 542898
rect 40794 507218 40826 507454
rect 41062 507218 41146 507454
rect 41382 507218 41414 507454
rect 40794 507134 41414 507218
rect 40794 506898 40826 507134
rect 41062 506898 41146 507134
rect 41382 506898 41414 507134
rect 40794 471454 41414 506898
rect 40794 471218 40826 471454
rect 41062 471218 41146 471454
rect 41382 471218 41414 471454
rect 40794 471134 41414 471218
rect 40794 470898 40826 471134
rect 41062 470898 41146 471134
rect 41382 470898 41414 471134
rect 40794 435454 41414 470898
rect 40794 435218 40826 435454
rect 41062 435218 41146 435454
rect 41382 435218 41414 435454
rect 40794 435134 41414 435218
rect 40794 434898 40826 435134
rect 41062 434898 41146 435134
rect 41382 434898 41414 435134
rect 40794 399454 41414 434898
rect 40794 399218 40826 399454
rect 41062 399218 41146 399454
rect 41382 399218 41414 399454
rect 40794 399134 41414 399218
rect 40794 398898 40826 399134
rect 41062 398898 41146 399134
rect 41382 398898 41414 399134
rect 40794 363454 41414 398898
rect 40794 363218 40826 363454
rect 41062 363218 41146 363454
rect 41382 363218 41414 363454
rect 40794 363134 41414 363218
rect 40794 362898 40826 363134
rect 41062 362898 41146 363134
rect 41382 362898 41414 363134
rect 40794 327454 41414 362898
rect 40794 327218 40826 327454
rect 41062 327218 41146 327454
rect 41382 327218 41414 327454
rect 40794 327134 41414 327218
rect 40794 326898 40826 327134
rect 41062 326898 41146 327134
rect 41382 326898 41414 327134
rect 40794 291454 41414 326898
rect 40794 291218 40826 291454
rect 41062 291218 41146 291454
rect 41382 291218 41414 291454
rect 40794 291134 41414 291218
rect 40794 290898 40826 291134
rect 41062 290898 41146 291134
rect 41382 290898 41414 291134
rect 40794 255454 41414 290898
rect 40794 255218 40826 255454
rect 41062 255218 41146 255454
rect 41382 255218 41414 255454
rect 40794 255134 41414 255218
rect 40794 254898 40826 255134
rect 41062 254898 41146 255134
rect 41382 254898 41414 255134
rect 40794 219454 41414 254898
rect 40794 219218 40826 219454
rect 41062 219218 41146 219454
rect 41382 219218 41414 219454
rect 40794 219134 41414 219218
rect 40794 218898 40826 219134
rect 41062 218898 41146 219134
rect 41382 218898 41414 219134
rect 40794 183454 41414 218898
rect 40794 183218 40826 183454
rect 41062 183218 41146 183454
rect 41382 183218 41414 183454
rect 40794 183134 41414 183218
rect 40794 182898 40826 183134
rect 41062 182898 41146 183134
rect 41382 182898 41414 183134
rect 40794 147454 41414 182898
rect 40794 147218 40826 147454
rect 41062 147218 41146 147454
rect 41382 147218 41414 147454
rect 40794 147134 41414 147218
rect 40794 146898 40826 147134
rect 41062 146898 41146 147134
rect 41382 146898 41414 147134
rect 40794 111454 41414 146898
rect 40794 111218 40826 111454
rect 41062 111218 41146 111454
rect 41382 111218 41414 111454
rect 40794 111134 41414 111218
rect 40794 110898 40826 111134
rect 41062 110898 41146 111134
rect 41382 110898 41414 111134
rect 40794 75454 41414 110898
rect 40794 75218 40826 75454
rect 41062 75218 41146 75454
rect 41382 75218 41414 75454
rect 40794 75134 41414 75218
rect 40794 74898 40826 75134
rect 41062 74898 41146 75134
rect 41382 74898 41414 75134
rect 40794 74295 41414 74898
rect 41954 680614 42574 711002
rect 51954 710598 52574 711590
rect 51954 710362 51986 710598
rect 52222 710362 52306 710598
rect 52542 710362 52574 710598
rect 51954 710278 52574 710362
rect 51954 710042 51986 710278
rect 52222 710042 52306 710278
rect 52542 710042 52574 710278
rect 48234 708678 48854 709670
rect 48234 708442 48266 708678
rect 48502 708442 48586 708678
rect 48822 708442 48854 708678
rect 48234 708358 48854 708442
rect 48234 708122 48266 708358
rect 48502 708122 48586 708358
rect 48822 708122 48854 708358
rect 41954 680378 41986 680614
rect 42222 680378 42306 680614
rect 42542 680378 42574 680614
rect 41954 680294 42574 680378
rect 41954 680058 41986 680294
rect 42222 680058 42306 680294
rect 42542 680058 42574 680294
rect 41954 644614 42574 680058
rect 41954 644378 41986 644614
rect 42222 644378 42306 644614
rect 42542 644378 42574 644614
rect 41954 644294 42574 644378
rect 41954 644058 41986 644294
rect 42222 644058 42306 644294
rect 42542 644058 42574 644294
rect 41954 608614 42574 644058
rect 41954 608378 41986 608614
rect 42222 608378 42306 608614
rect 42542 608378 42574 608614
rect 41954 608294 42574 608378
rect 41954 608058 41986 608294
rect 42222 608058 42306 608294
rect 42542 608058 42574 608294
rect 41954 572614 42574 608058
rect 41954 572378 41986 572614
rect 42222 572378 42306 572614
rect 42542 572378 42574 572614
rect 41954 572294 42574 572378
rect 41954 572058 41986 572294
rect 42222 572058 42306 572294
rect 42542 572058 42574 572294
rect 41954 536614 42574 572058
rect 41954 536378 41986 536614
rect 42222 536378 42306 536614
rect 42542 536378 42574 536614
rect 41954 536294 42574 536378
rect 41954 536058 41986 536294
rect 42222 536058 42306 536294
rect 42542 536058 42574 536294
rect 41954 500614 42574 536058
rect 41954 500378 41986 500614
rect 42222 500378 42306 500614
rect 42542 500378 42574 500614
rect 41954 500294 42574 500378
rect 41954 500058 41986 500294
rect 42222 500058 42306 500294
rect 42542 500058 42574 500294
rect 41954 464614 42574 500058
rect 41954 464378 41986 464614
rect 42222 464378 42306 464614
rect 42542 464378 42574 464614
rect 41954 464294 42574 464378
rect 41954 464058 41986 464294
rect 42222 464058 42306 464294
rect 42542 464058 42574 464294
rect 41954 428614 42574 464058
rect 41954 428378 41986 428614
rect 42222 428378 42306 428614
rect 42542 428378 42574 428614
rect 41954 428294 42574 428378
rect 41954 428058 41986 428294
rect 42222 428058 42306 428294
rect 42542 428058 42574 428294
rect 41954 392614 42574 428058
rect 41954 392378 41986 392614
rect 42222 392378 42306 392614
rect 42542 392378 42574 392614
rect 41954 392294 42574 392378
rect 41954 392058 41986 392294
rect 42222 392058 42306 392294
rect 42542 392058 42574 392294
rect 41954 356614 42574 392058
rect 41954 356378 41986 356614
rect 42222 356378 42306 356614
rect 42542 356378 42574 356614
rect 41954 356294 42574 356378
rect 41954 356058 41986 356294
rect 42222 356058 42306 356294
rect 42542 356058 42574 356294
rect 41954 320614 42574 356058
rect 41954 320378 41986 320614
rect 42222 320378 42306 320614
rect 42542 320378 42574 320614
rect 41954 320294 42574 320378
rect 41954 320058 41986 320294
rect 42222 320058 42306 320294
rect 42542 320058 42574 320294
rect 41954 284614 42574 320058
rect 41954 284378 41986 284614
rect 42222 284378 42306 284614
rect 42542 284378 42574 284614
rect 41954 284294 42574 284378
rect 41954 284058 41986 284294
rect 42222 284058 42306 284294
rect 42542 284058 42574 284294
rect 41954 248614 42574 284058
rect 41954 248378 41986 248614
rect 42222 248378 42306 248614
rect 42542 248378 42574 248614
rect 41954 248294 42574 248378
rect 41954 248058 41986 248294
rect 42222 248058 42306 248294
rect 42542 248058 42574 248294
rect 41954 212614 42574 248058
rect 41954 212378 41986 212614
rect 42222 212378 42306 212614
rect 42542 212378 42574 212614
rect 41954 212294 42574 212378
rect 41954 212058 41986 212294
rect 42222 212058 42306 212294
rect 42542 212058 42574 212294
rect 41954 176614 42574 212058
rect 41954 176378 41986 176614
rect 42222 176378 42306 176614
rect 42542 176378 42574 176614
rect 41954 176294 42574 176378
rect 41954 176058 41986 176294
rect 42222 176058 42306 176294
rect 42542 176058 42574 176294
rect 41954 140614 42574 176058
rect 41954 140378 41986 140614
rect 42222 140378 42306 140614
rect 42542 140378 42574 140614
rect 41954 140294 42574 140378
rect 41954 140058 41986 140294
rect 42222 140058 42306 140294
rect 42542 140058 42574 140294
rect 41954 104614 42574 140058
rect 41954 104378 41986 104614
rect 42222 104378 42306 104614
rect 42542 104378 42574 104614
rect 41954 104294 42574 104378
rect 41954 104058 41986 104294
rect 42222 104058 42306 104294
rect 42542 104058 42574 104294
rect 41954 74295 42574 104058
rect 44514 706758 45134 707750
rect 44514 706522 44546 706758
rect 44782 706522 44866 706758
rect 45102 706522 45134 706758
rect 44514 706438 45134 706522
rect 44514 706202 44546 706438
rect 44782 706202 44866 706438
rect 45102 706202 45134 706438
rect 44514 691174 45134 706202
rect 44514 690938 44546 691174
rect 44782 690938 44866 691174
rect 45102 690938 45134 691174
rect 44514 690854 45134 690938
rect 44514 690618 44546 690854
rect 44782 690618 44866 690854
rect 45102 690618 45134 690854
rect 44514 655174 45134 690618
rect 44514 654938 44546 655174
rect 44782 654938 44866 655174
rect 45102 654938 45134 655174
rect 44514 654854 45134 654938
rect 44514 654618 44546 654854
rect 44782 654618 44866 654854
rect 45102 654618 45134 654854
rect 44514 619174 45134 654618
rect 44514 618938 44546 619174
rect 44782 618938 44866 619174
rect 45102 618938 45134 619174
rect 44514 618854 45134 618938
rect 44514 618618 44546 618854
rect 44782 618618 44866 618854
rect 45102 618618 45134 618854
rect 44514 583174 45134 618618
rect 44514 582938 44546 583174
rect 44782 582938 44866 583174
rect 45102 582938 45134 583174
rect 44514 582854 45134 582938
rect 44514 582618 44546 582854
rect 44782 582618 44866 582854
rect 45102 582618 45134 582854
rect 44514 547174 45134 582618
rect 44514 546938 44546 547174
rect 44782 546938 44866 547174
rect 45102 546938 45134 547174
rect 44514 546854 45134 546938
rect 44514 546618 44546 546854
rect 44782 546618 44866 546854
rect 45102 546618 45134 546854
rect 44514 511174 45134 546618
rect 44514 510938 44546 511174
rect 44782 510938 44866 511174
rect 45102 510938 45134 511174
rect 44514 510854 45134 510938
rect 44514 510618 44546 510854
rect 44782 510618 44866 510854
rect 45102 510618 45134 510854
rect 44514 475174 45134 510618
rect 44514 474938 44546 475174
rect 44782 474938 44866 475174
rect 45102 474938 45134 475174
rect 44514 474854 45134 474938
rect 44514 474618 44546 474854
rect 44782 474618 44866 474854
rect 45102 474618 45134 474854
rect 44514 439174 45134 474618
rect 44514 438938 44546 439174
rect 44782 438938 44866 439174
rect 45102 438938 45134 439174
rect 44514 438854 45134 438938
rect 44514 438618 44546 438854
rect 44782 438618 44866 438854
rect 45102 438618 45134 438854
rect 44514 403174 45134 438618
rect 44514 402938 44546 403174
rect 44782 402938 44866 403174
rect 45102 402938 45134 403174
rect 44514 402854 45134 402938
rect 44514 402618 44546 402854
rect 44782 402618 44866 402854
rect 45102 402618 45134 402854
rect 44514 367174 45134 402618
rect 44514 366938 44546 367174
rect 44782 366938 44866 367174
rect 45102 366938 45134 367174
rect 44514 366854 45134 366938
rect 44514 366618 44546 366854
rect 44782 366618 44866 366854
rect 45102 366618 45134 366854
rect 44514 331174 45134 366618
rect 44514 330938 44546 331174
rect 44782 330938 44866 331174
rect 45102 330938 45134 331174
rect 44514 330854 45134 330938
rect 44514 330618 44546 330854
rect 44782 330618 44866 330854
rect 45102 330618 45134 330854
rect 44514 295174 45134 330618
rect 44514 294938 44546 295174
rect 44782 294938 44866 295174
rect 45102 294938 45134 295174
rect 44514 294854 45134 294938
rect 44514 294618 44546 294854
rect 44782 294618 44866 294854
rect 45102 294618 45134 294854
rect 44514 259174 45134 294618
rect 44514 258938 44546 259174
rect 44782 258938 44866 259174
rect 45102 258938 45134 259174
rect 44514 258854 45134 258938
rect 44514 258618 44546 258854
rect 44782 258618 44866 258854
rect 45102 258618 45134 258854
rect 44514 223174 45134 258618
rect 44514 222938 44546 223174
rect 44782 222938 44866 223174
rect 45102 222938 45134 223174
rect 44514 222854 45134 222938
rect 44514 222618 44546 222854
rect 44782 222618 44866 222854
rect 45102 222618 45134 222854
rect 44514 187174 45134 222618
rect 44514 186938 44546 187174
rect 44782 186938 44866 187174
rect 45102 186938 45134 187174
rect 44514 186854 45134 186938
rect 44514 186618 44546 186854
rect 44782 186618 44866 186854
rect 45102 186618 45134 186854
rect 44514 151174 45134 186618
rect 44514 150938 44546 151174
rect 44782 150938 44866 151174
rect 45102 150938 45134 151174
rect 44514 150854 45134 150938
rect 44514 150618 44546 150854
rect 44782 150618 44866 150854
rect 45102 150618 45134 150854
rect 44514 115174 45134 150618
rect 44514 114938 44546 115174
rect 44782 114938 44866 115174
rect 45102 114938 45134 115174
rect 44514 114854 45134 114938
rect 44514 114618 44546 114854
rect 44782 114618 44866 114854
rect 45102 114618 45134 114854
rect 44514 79174 45134 114618
rect 44514 78938 44546 79174
rect 44782 78938 44866 79174
rect 45102 78938 45134 79174
rect 44514 78854 45134 78938
rect 44514 78618 44546 78854
rect 44782 78618 44866 78854
rect 45102 78618 45134 78854
rect 44514 74295 45134 78618
rect 48234 694894 48854 708122
rect 48234 694658 48266 694894
rect 48502 694658 48586 694894
rect 48822 694658 48854 694894
rect 48234 694574 48854 694658
rect 48234 694338 48266 694574
rect 48502 694338 48586 694574
rect 48822 694338 48854 694574
rect 48234 658894 48854 694338
rect 48234 658658 48266 658894
rect 48502 658658 48586 658894
rect 48822 658658 48854 658894
rect 48234 658574 48854 658658
rect 48234 658338 48266 658574
rect 48502 658338 48586 658574
rect 48822 658338 48854 658574
rect 48234 622894 48854 658338
rect 48234 622658 48266 622894
rect 48502 622658 48586 622894
rect 48822 622658 48854 622894
rect 48234 622574 48854 622658
rect 48234 622338 48266 622574
rect 48502 622338 48586 622574
rect 48822 622338 48854 622574
rect 48234 586894 48854 622338
rect 48234 586658 48266 586894
rect 48502 586658 48586 586894
rect 48822 586658 48854 586894
rect 48234 586574 48854 586658
rect 48234 586338 48266 586574
rect 48502 586338 48586 586574
rect 48822 586338 48854 586574
rect 48234 550894 48854 586338
rect 48234 550658 48266 550894
rect 48502 550658 48586 550894
rect 48822 550658 48854 550894
rect 48234 550574 48854 550658
rect 48234 550338 48266 550574
rect 48502 550338 48586 550574
rect 48822 550338 48854 550574
rect 48234 514894 48854 550338
rect 48234 514658 48266 514894
rect 48502 514658 48586 514894
rect 48822 514658 48854 514894
rect 48234 514574 48854 514658
rect 48234 514338 48266 514574
rect 48502 514338 48586 514574
rect 48822 514338 48854 514574
rect 48234 478894 48854 514338
rect 48234 478658 48266 478894
rect 48502 478658 48586 478894
rect 48822 478658 48854 478894
rect 48234 478574 48854 478658
rect 48234 478338 48266 478574
rect 48502 478338 48586 478574
rect 48822 478338 48854 478574
rect 48234 442894 48854 478338
rect 48234 442658 48266 442894
rect 48502 442658 48586 442894
rect 48822 442658 48854 442894
rect 48234 442574 48854 442658
rect 48234 442338 48266 442574
rect 48502 442338 48586 442574
rect 48822 442338 48854 442574
rect 48234 406894 48854 442338
rect 48234 406658 48266 406894
rect 48502 406658 48586 406894
rect 48822 406658 48854 406894
rect 48234 406574 48854 406658
rect 48234 406338 48266 406574
rect 48502 406338 48586 406574
rect 48822 406338 48854 406574
rect 48234 370894 48854 406338
rect 48234 370658 48266 370894
rect 48502 370658 48586 370894
rect 48822 370658 48854 370894
rect 48234 370574 48854 370658
rect 48234 370338 48266 370574
rect 48502 370338 48586 370574
rect 48822 370338 48854 370574
rect 48234 334894 48854 370338
rect 48234 334658 48266 334894
rect 48502 334658 48586 334894
rect 48822 334658 48854 334894
rect 48234 334574 48854 334658
rect 48234 334338 48266 334574
rect 48502 334338 48586 334574
rect 48822 334338 48854 334574
rect 48234 298894 48854 334338
rect 48234 298658 48266 298894
rect 48502 298658 48586 298894
rect 48822 298658 48854 298894
rect 48234 298574 48854 298658
rect 48234 298338 48266 298574
rect 48502 298338 48586 298574
rect 48822 298338 48854 298574
rect 48234 262894 48854 298338
rect 48234 262658 48266 262894
rect 48502 262658 48586 262894
rect 48822 262658 48854 262894
rect 48234 262574 48854 262658
rect 48234 262338 48266 262574
rect 48502 262338 48586 262574
rect 48822 262338 48854 262574
rect 48234 226894 48854 262338
rect 48234 226658 48266 226894
rect 48502 226658 48586 226894
rect 48822 226658 48854 226894
rect 48234 226574 48854 226658
rect 48234 226338 48266 226574
rect 48502 226338 48586 226574
rect 48822 226338 48854 226574
rect 48234 190894 48854 226338
rect 48234 190658 48266 190894
rect 48502 190658 48586 190894
rect 48822 190658 48854 190894
rect 48234 190574 48854 190658
rect 48234 190338 48266 190574
rect 48502 190338 48586 190574
rect 48822 190338 48854 190574
rect 48234 154894 48854 190338
rect 48234 154658 48266 154894
rect 48502 154658 48586 154894
rect 48822 154658 48854 154894
rect 48234 154574 48854 154658
rect 48234 154338 48266 154574
rect 48502 154338 48586 154574
rect 48822 154338 48854 154574
rect 48234 118894 48854 154338
rect 48234 118658 48266 118894
rect 48502 118658 48586 118894
rect 48822 118658 48854 118894
rect 48234 118574 48854 118658
rect 48234 118338 48266 118574
rect 48502 118338 48586 118574
rect 48822 118338 48854 118574
rect 48234 82894 48854 118338
rect 48234 82658 48266 82894
rect 48502 82658 48586 82894
rect 48822 82658 48854 82894
rect 48234 82574 48854 82658
rect 48234 82338 48266 82574
rect 48502 82338 48586 82574
rect 48822 82338 48854 82574
rect 48234 74295 48854 82338
rect 50794 705798 51414 705830
rect 50794 705562 50826 705798
rect 51062 705562 51146 705798
rect 51382 705562 51414 705798
rect 50794 705478 51414 705562
rect 50794 705242 50826 705478
rect 51062 705242 51146 705478
rect 51382 705242 51414 705478
rect 50794 669454 51414 705242
rect 50794 669218 50826 669454
rect 51062 669218 51146 669454
rect 51382 669218 51414 669454
rect 50794 669134 51414 669218
rect 50794 668898 50826 669134
rect 51062 668898 51146 669134
rect 51382 668898 51414 669134
rect 50794 633454 51414 668898
rect 50794 633218 50826 633454
rect 51062 633218 51146 633454
rect 51382 633218 51414 633454
rect 50794 633134 51414 633218
rect 50794 632898 50826 633134
rect 51062 632898 51146 633134
rect 51382 632898 51414 633134
rect 50794 597454 51414 632898
rect 50794 597218 50826 597454
rect 51062 597218 51146 597454
rect 51382 597218 51414 597454
rect 50794 597134 51414 597218
rect 50794 596898 50826 597134
rect 51062 596898 51146 597134
rect 51382 596898 51414 597134
rect 50794 561454 51414 596898
rect 50794 561218 50826 561454
rect 51062 561218 51146 561454
rect 51382 561218 51414 561454
rect 50794 561134 51414 561218
rect 50794 560898 50826 561134
rect 51062 560898 51146 561134
rect 51382 560898 51414 561134
rect 50794 525454 51414 560898
rect 50794 525218 50826 525454
rect 51062 525218 51146 525454
rect 51382 525218 51414 525454
rect 50794 525134 51414 525218
rect 50794 524898 50826 525134
rect 51062 524898 51146 525134
rect 51382 524898 51414 525134
rect 50794 489454 51414 524898
rect 50794 489218 50826 489454
rect 51062 489218 51146 489454
rect 51382 489218 51414 489454
rect 50794 489134 51414 489218
rect 50794 488898 50826 489134
rect 51062 488898 51146 489134
rect 51382 488898 51414 489134
rect 50794 453454 51414 488898
rect 50794 453218 50826 453454
rect 51062 453218 51146 453454
rect 51382 453218 51414 453454
rect 50794 453134 51414 453218
rect 50794 452898 50826 453134
rect 51062 452898 51146 453134
rect 51382 452898 51414 453134
rect 50794 417454 51414 452898
rect 50794 417218 50826 417454
rect 51062 417218 51146 417454
rect 51382 417218 51414 417454
rect 50794 417134 51414 417218
rect 50794 416898 50826 417134
rect 51062 416898 51146 417134
rect 51382 416898 51414 417134
rect 50794 381454 51414 416898
rect 50794 381218 50826 381454
rect 51062 381218 51146 381454
rect 51382 381218 51414 381454
rect 50794 381134 51414 381218
rect 50794 380898 50826 381134
rect 51062 380898 51146 381134
rect 51382 380898 51414 381134
rect 50794 345454 51414 380898
rect 50794 345218 50826 345454
rect 51062 345218 51146 345454
rect 51382 345218 51414 345454
rect 50794 345134 51414 345218
rect 50794 344898 50826 345134
rect 51062 344898 51146 345134
rect 51382 344898 51414 345134
rect 50794 309454 51414 344898
rect 50794 309218 50826 309454
rect 51062 309218 51146 309454
rect 51382 309218 51414 309454
rect 50794 309134 51414 309218
rect 50794 308898 50826 309134
rect 51062 308898 51146 309134
rect 51382 308898 51414 309134
rect 50794 273454 51414 308898
rect 50794 273218 50826 273454
rect 51062 273218 51146 273454
rect 51382 273218 51414 273454
rect 50794 273134 51414 273218
rect 50794 272898 50826 273134
rect 51062 272898 51146 273134
rect 51382 272898 51414 273134
rect 50794 237454 51414 272898
rect 50794 237218 50826 237454
rect 51062 237218 51146 237454
rect 51382 237218 51414 237454
rect 50794 237134 51414 237218
rect 50794 236898 50826 237134
rect 51062 236898 51146 237134
rect 51382 236898 51414 237134
rect 50794 201454 51414 236898
rect 50794 201218 50826 201454
rect 51062 201218 51146 201454
rect 51382 201218 51414 201454
rect 50794 201134 51414 201218
rect 50794 200898 50826 201134
rect 51062 200898 51146 201134
rect 51382 200898 51414 201134
rect 50794 165454 51414 200898
rect 50794 165218 50826 165454
rect 51062 165218 51146 165454
rect 51382 165218 51414 165454
rect 50794 165134 51414 165218
rect 50794 164898 50826 165134
rect 51062 164898 51146 165134
rect 51382 164898 51414 165134
rect 50794 129454 51414 164898
rect 50794 129218 50826 129454
rect 51062 129218 51146 129454
rect 51382 129218 51414 129454
rect 50794 129134 51414 129218
rect 50794 128898 50826 129134
rect 51062 128898 51146 129134
rect 51382 128898 51414 129134
rect 50794 93454 51414 128898
rect 50794 93218 50826 93454
rect 51062 93218 51146 93454
rect 51382 93218 51414 93454
rect 50794 93134 51414 93218
rect 50794 92898 50826 93134
rect 51062 92898 51146 93134
rect 51382 92898 51414 93134
rect 50794 74295 51414 92898
rect 51954 698614 52574 710042
rect 61954 711558 62574 711590
rect 61954 711322 61986 711558
rect 62222 711322 62306 711558
rect 62542 711322 62574 711558
rect 61954 711238 62574 711322
rect 61954 711002 61986 711238
rect 62222 711002 62306 711238
rect 62542 711002 62574 711238
rect 58234 709638 58854 709670
rect 58234 709402 58266 709638
rect 58502 709402 58586 709638
rect 58822 709402 58854 709638
rect 58234 709318 58854 709402
rect 58234 709082 58266 709318
rect 58502 709082 58586 709318
rect 58822 709082 58854 709318
rect 51954 698378 51986 698614
rect 52222 698378 52306 698614
rect 52542 698378 52574 698614
rect 51954 698294 52574 698378
rect 51954 698058 51986 698294
rect 52222 698058 52306 698294
rect 52542 698058 52574 698294
rect 51954 662614 52574 698058
rect 51954 662378 51986 662614
rect 52222 662378 52306 662614
rect 52542 662378 52574 662614
rect 51954 662294 52574 662378
rect 51954 662058 51986 662294
rect 52222 662058 52306 662294
rect 52542 662058 52574 662294
rect 51954 626614 52574 662058
rect 51954 626378 51986 626614
rect 52222 626378 52306 626614
rect 52542 626378 52574 626614
rect 51954 626294 52574 626378
rect 51954 626058 51986 626294
rect 52222 626058 52306 626294
rect 52542 626058 52574 626294
rect 51954 590614 52574 626058
rect 51954 590378 51986 590614
rect 52222 590378 52306 590614
rect 52542 590378 52574 590614
rect 51954 590294 52574 590378
rect 51954 590058 51986 590294
rect 52222 590058 52306 590294
rect 52542 590058 52574 590294
rect 51954 554614 52574 590058
rect 51954 554378 51986 554614
rect 52222 554378 52306 554614
rect 52542 554378 52574 554614
rect 51954 554294 52574 554378
rect 51954 554058 51986 554294
rect 52222 554058 52306 554294
rect 52542 554058 52574 554294
rect 51954 518614 52574 554058
rect 51954 518378 51986 518614
rect 52222 518378 52306 518614
rect 52542 518378 52574 518614
rect 51954 518294 52574 518378
rect 51954 518058 51986 518294
rect 52222 518058 52306 518294
rect 52542 518058 52574 518294
rect 51954 482614 52574 518058
rect 51954 482378 51986 482614
rect 52222 482378 52306 482614
rect 52542 482378 52574 482614
rect 51954 482294 52574 482378
rect 51954 482058 51986 482294
rect 52222 482058 52306 482294
rect 52542 482058 52574 482294
rect 51954 446614 52574 482058
rect 51954 446378 51986 446614
rect 52222 446378 52306 446614
rect 52542 446378 52574 446614
rect 51954 446294 52574 446378
rect 51954 446058 51986 446294
rect 52222 446058 52306 446294
rect 52542 446058 52574 446294
rect 51954 410614 52574 446058
rect 51954 410378 51986 410614
rect 52222 410378 52306 410614
rect 52542 410378 52574 410614
rect 51954 410294 52574 410378
rect 51954 410058 51986 410294
rect 52222 410058 52306 410294
rect 52542 410058 52574 410294
rect 51954 374614 52574 410058
rect 51954 374378 51986 374614
rect 52222 374378 52306 374614
rect 52542 374378 52574 374614
rect 51954 374294 52574 374378
rect 51954 374058 51986 374294
rect 52222 374058 52306 374294
rect 52542 374058 52574 374294
rect 51954 338614 52574 374058
rect 51954 338378 51986 338614
rect 52222 338378 52306 338614
rect 52542 338378 52574 338614
rect 51954 338294 52574 338378
rect 51954 338058 51986 338294
rect 52222 338058 52306 338294
rect 52542 338058 52574 338294
rect 51954 302614 52574 338058
rect 51954 302378 51986 302614
rect 52222 302378 52306 302614
rect 52542 302378 52574 302614
rect 51954 302294 52574 302378
rect 51954 302058 51986 302294
rect 52222 302058 52306 302294
rect 52542 302058 52574 302294
rect 51954 266614 52574 302058
rect 51954 266378 51986 266614
rect 52222 266378 52306 266614
rect 52542 266378 52574 266614
rect 51954 266294 52574 266378
rect 51954 266058 51986 266294
rect 52222 266058 52306 266294
rect 52542 266058 52574 266294
rect 51954 230614 52574 266058
rect 51954 230378 51986 230614
rect 52222 230378 52306 230614
rect 52542 230378 52574 230614
rect 51954 230294 52574 230378
rect 51954 230058 51986 230294
rect 52222 230058 52306 230294
rect 52542 230058 52574 230294
rect 51954 194614 52574 230058
rect 51954 194378 51986 194614
rect 52222 194378 52306 194614
rect 52542 194378 52574 194614
rect 51954 194294 52574 194378
rect 51954 194058 51986 194294
rect 52222 194058 52306 194294
rect 52542 194058 52574 194294
rect 51954 158614 52574 194058
rect 51954 158378 51986 158614
rect 52222 158378 52306 158614
rect 52542 158378 52574 158614
rect 51954 158294 52574 158378
rect 51954 158058 51986 158294
rect 52222 158058 52306 158294
rect 52542 158058 52574 158294
rect 51954 122614 52574 158058
rect 51954 122378 51986 122614
rect 52222 122378 52306 122614
rect 52542 122378 52574 122614
rect 51954 122294 52574 122378
rect 51954 122058 51986 122294
rect 52222 122058 52306 122294
rect 52542 122058 52574 122294
rect 51954 86614 52574 122058
rect 51954 86378 51986 86614
rect 52222 86378 52306 86614
rect 52542 86378 52574 86614
rect 51954 86294 52574 86378
rect 51954 86058 51986 86294
rect 52222 86058 52306 86294
rect 52542 86058 52574 86294
rect 51954 74295 52574 86058
rect 54514 707718 55134 707750
rect 54514 707482 54546 707718
rect 54782 707482 54866 707718
rect 55102 707482 55134 707718
rect 54514 707398 55134 707482
rect 54514 707162 54546 707398
rect 54782 707162 54866 707398
rect 55102 707162 55134 707398
rect 54514 673174 55134 707162
rect 54514 672938 54546 673174
rect 54782 672938 54866 673174
rect 55102 672938 55134 673174
rect 54514 672854 55134 672938
rect 54514 672618 54546 672854
rect 54782 672618 54866 672854
rect 55102 672618 55134 672854
rect 54514 637174 55134 672618
rect 54514 636938 54546 637174
rect 54782 636938 54866 637174
rect 55102 636938 55134 637174
rect 54514 636854 55134 636938
rect 54514 636618 54546 636854
rect 54782 636618 54866 636854
rect 55102 636618 55134 636854
rect 54514 601174 55134 636618
rect 54514 600938 54546 601174
rect 54782 600938 54866 601174
rect 55102 600938 55134 601174
rect 54514 600854 55134 600938
rect 54514 600618 54546 600854
rect 54782 600618 54866 600854
rect 55102 600618 55134 600854
rect 54514 565174 55134 600618
rect 54514 564938 54546 565174
rect 54782 564938 54866 565174
rect 55102 564938 55134 565174
rect 54514 564854 55134 564938
rect 54514 564618 54546 564854
rect 54782 564618 54866 564854
rect 55102 564618 55134 564854
rect 54514 529174 55134 564618
rect 54514 528938 54546 529174
rect 54782 528938 54866 529174
rect 55102 528938 55134 529174
rect 54514 528854 55134 528938
rect 54514 528618 54546 528854
rect 54782 528618 54866 528854
rect 55102 528618 55134 528854
rect 54514 493174 55134 528618
rect 54514 492938 54546 493174
rect 54782 492938 54866 493174
rect 55102 492938 55134 493174
rect 54514 492854 55134 492938
rect 54514 492618 54546 492854
rect 54782 492618 54866 492854
rect 55102 492618 55134 492854
rect 54514 457174 55134 492618
rect 54514 456938 54546 457174
rect 54782 456938 54866 457174
rect 55102 456938 55134 457174
rect 54514 456854 55134 456938
rect 54514 456618 54546 456854
rect 54782 456618 54866 456854
rect 55102 456618 55134 456854
rect 54514 421174 55134 456618
rect 54514 420938 54546 421174
rect 54782 420938 54866 421174
rect 55102 420938 55134 421174
rect 54514 420854 55134 420938
rect 54514 420618 54546 420854
rect 54782 420618 54866 420854
rect 55102 420618 55134 420854
rect 54514 385174 55134 420618
rect 54514 384938 54546 385174
rect 54782 384938 54866 385174
rect 55102 384938 55134 385174
rect 54514 384854 55134 384938
rect 54514 384618 54546 384854
rect 54782 384618 54866 384854
rect 55102 384618 55134 384854
rect 54514 349174 55134 384618
rect 54514 348938 54546 349174
rect 54782 348938 54866 349174
rect 55102 348938 55134 349174
rect 54514 348854 55134 348938
rect 54514 348618 54546 348854
rect 54782 348618 54866 348854
rect 55102 348618 55134 348854
rect 54514 313174 55134 348618
rect 54514 312938 54546 313174
rect 54782 312938 54866 313174
rect 55102 312938 55134 313174
rect 54514 312854 55134 312938
rect 54514 312618 54546 312854
rect 54782 312618 54866 312854
rect 55102 312618 55134 312854
rect 54514 277174 55134 312618
rect 54514 276938 54546 277174
rect 54782 276938 54866 277174
rect 55102 276938 55134 277174
rect 54514 276854 55134 276938
rect 54514 276618 54546 276854
rect 54782 276618 54866 276854
rect 55102 276618 55134 276854
rect 54514 241174 55134 276618
rect 54514 240938 54546 241174
rect 54782 240938 54866 241174
rect 55102 240938 55134 241174
rect 54514 240854 55134 240938
rect 54514 240618 54546 240854
rect 54782 240618 54866 240854
rect 55102 240618 55134 240854
rect 54514 205174 55134 240618
rect 54514 204938 54546 205174
rect 54782 204938 54866 205174
rect 55102 204938 55134 205174
rect 54514 204854 55134 204938
rect 54514 204618 54546 204854
rect 54782 204618 54866 204854
rect 55102 204618 55134 204854
rect 54514 169174 55134 204618
rect 54514 168938 54546 169174
rect 54782 168938 54866 169174
rect 55102 168938 55134 169174
rect 54514 168854 55134 168938
rect 54514 168618 54546 168854
rect 54782 168618 54866 168854
rect 55102 168618 55134 168854
rect 54514 133174 55134 168618
rect 54514 132938 54546 133174
rect 54782 132938 54866 133174
rect 55102 132938 55134 133174
rect 54514 132854 55134 132938
rect 54514 132618 54546 132854
rect 54782 132618 54866 132854
rect 55102 132618 55134 132854
rect 54514 97174 55134 132618
rect 54514 96938 54546 97174
rect 54782 96938 54866 97174
rect 55102 96938 55134 97174
rect 54514 96854 55134 96938
rect 54514 96618 54546 96854
rect 54782 96618 54866 96854
rect 55102 96618 55134 96854
rect 54514 74295 55134 96618
rect 58234 676894 58854 709082
rect 58234 676658 58266 676894
rect 58502 676658 58586 676894
rect 58822 676658 58854 676894
rect 58234 676574 58854 676658
rect 58234 676338 58266 676574
rect 58502 676338 58586 676574
rect 58822 676338 58854 676574
rect 58234 640894 58854 676338
rect 58234 640658 58266 640894
rect 58502 640658 58586 640894
rect 58822 640658 58854 640894
rect 58234 640574 58854 640658
rect 58234 640338 58266 640574
rect 58502 640338 58586 640574
rect 58822 640338 58854 640574
rect 58234 604894 58854 640338
rect 58234 604658 58266 604894
rect 58502 604658 58586 604894
rect 58822 604658 58854 604894
rect 58234 604574 58854 604658
rect 58234 604338 58266 604574
rect 58502 604338 58586 604574
rect 58822 604338 58854 604574
rect 58234 568894 58854 604338
rect 58234 568658 58266 568894
rect 58502 568658 58586 568894
rect 58822 568658 58854 568894
rect 58234 568574 58854 568658
rect 58234 568338 58266 568574
rect 58502 568338 58586 568574
rect 58822 568338 58854 568574
rect 58234 532894 58854 568338
rect 58234 532658 58266 532894
rect 58502 532658 58586 532894
rect 58822 532658 58854 532894
rect 58234 532574 58854 532658
rect 58234 532338 58266 532574
rect 58502 532338 58586 532574
rect 58822 532338 58854 532574
rect 58234 496894 58854 532338
rect 58234 496658 58266 496894
rect 58502 496658 58586 496894
rect 58822 496658 58854 496894
rect 58234 496574 58854 496658
rect 58234 496338 58266 496574
rect 58502 496338 58586 496574
rect 58822 496338 58854 496574
rect 58234 460894 58854 496338
rect 58234 460658 58266 460894
rect 58502 460658 58586 460894
rect 58822 460658 58854 460894
rect 58234 460574 58854 460658
rect 58234 460338 58266 460574
rect 58502 460338 58586 460574
rect 58822 460338 58854 460574
rect 58234 424894 58854 460338
rect 58234 424658 58266 424894
rect 58502 424658 58586 424894
rect 58822 424658 58854 424894
rect 58234 424574 58854 424658
rect 58234 424338 58266 424574
rect 58502 424338 58586 424574
rect 58822 424338 58854 424574
rect 58234 388894 58854 424338
rect 58234 388658 58266 388894
rect 58502 388658 58586 388894
rect 58822 388658 58854 388894
rect 58234 388574 58854 388658
rect 58234 388338 58266 388574
rect 58502 388338 58586 388574
rect 58822 388338 58854 388574
rect 58234 352894 58854 388338
rect 58234 352658 58266 352894
rect 58502 352658 58586 352894
rect 58822 352658 58854 352894
rect 58234 352574 58854 352658
rect 58234 352338 58266 352574
rect 58502 352338 58586 352574
rect 58822 352338 58854 352574
rect 58234 316894 58854 352338
rect 58234 316658 58266 316894
rect 58502 316658 58586 316894
rect 58822 316658 58854 316894
rect 58234 316574 58854 316658
rect 58234 316338 58266 316574
rect 58502 316338 58586 316574
rect 58822 316338 58854 316574
rect 58234 280894 58854 316338
rect 58234 280658 58266 280894
rect 58502 280658 58586 280894
rect 58822 280658 58854 280894
rect 58234 280574 58854 280658
rect 58234 280338 58266 280574
rect 58502 280338 58586 280574
rect 58822 280338 58854 280574
rect 58234 244894 58854 280338
rect 58234 244658 58266 244894
rect 58502 244658 58586 244894
rect 58822 244658 58854 244894
rect 58234 244574 58854 244658
rect 58234 244338 58266 244574
rect 58502 244338 58586 244574
rect 58822 244338 58854 244574
rect 58234 208894 58854 244338
rect 58234 208658 58266 208894
rect 58502 208658 58586 208894
rect 58822 208658 58854 208894
rect 58234 208574 58854 208658
rect 58234 208338 58266 208574
rect 58502 208338 58586 208574
rect 58822 208338 58854 208574
rect 58234 172894 58854 208338
rect 58234 172658 58266 172894
rect 58502 172658 58586 172894
rect 58822 172658 58854 172894
rect 58234 172574 58854 172658
rect 58234 172338 58266 172574
rect 58502 172338 58586 172574
rect 58822 172338 58854 172574
rect 58234 136894 58854 172338
rect 58234 136658 58266 136894
rect 58502 136658 58586 136894
rect 58822 136658 58854 136894
rect 58234 136574 58854 136658
rect 58234 136338 58266 136574
rect 58502 136338 58586 136574
rect 58822 136338 58854 136574
rect 58234 100894 58854 136338
rect 58234 100658 58266 100894
rect 58502 100658 58586 100894
rect 58822 100658 58854 100894
rect 58234 100574 58854 100658
rect 58234 100338 58266 100574
rect 58502 100338 58586 100574
rect 58822 100338 58854 100574
rect 58234 74295 58854 100338
rect 60794 704838 61414 705830
rect 60794 704602 60826 704838
rect 61062 704602 61146 704838
rect 61382 704602 61414 704838
rect 60794 704518 61414 704602
rect 60794 704282 60826 704518
rect 61062 704282 61146 704518
rect 61382 704282 61414 704518
rect 60794 687454 61414 704282
rect 60794 687218 60826 687454
rect 61062 687218 61146 687454
rect 61382 687218 61414 687454
rect 60794 687134 61414 687218
rect 60794 686898 60826 687134
rect 61062 686898 61146 687134
rect 61382 686898 61414 687134
rect 60794 651454 61414 686898
rect 60794 651218 60826 651454
rect 61062 651218 61146 651454
rect 61382 651218 61414 651454
rect 60794 651134 61414 651218
rect 60794 650898 60826 651134
rect 61062 650898 61146 651134
rect 61382 650898 61414 651134
rect 60794 615454 61414 650898
rect 60794 615218 60826 615454
rect 61062 615218 61146 615454
rect 61382 615218 61414 615454
rect 60794 615134 61414 615218
rect 60794 614898 60826 615134
rect 61062 614898 61146 615134
rect 61382 614898 61414 615134
rect 60794 579454 61414 614898
rect 60794 579218 60826 579454
rect 61062 579218 61146 579454
rect 61382 579218 61414 579454
rect 60794 579134 61414 579218
rect 60794 578898 60826 579134
rect 61062 578898 61146 579134
rect 61382 578898 61414 579134
rect 60794 543454 61414 578898
rect 60794 543218 60826 543454
rect 61062 543218 61146 543454
rect 61382 543218 61414 543454
rect 60794 543134 61414 543218
rect 60794 542898 60826 543134
rect 61062 542898 61146 543134
rect 61382 542898 61414 543134
rect 60794 507454 61414 542898
rect 60794 507218 60826 507454
rect 61062 507218 61146 507454
rect 61382 507218 61414 507454
rect 60794 507134 61414 507218
rect 60794 506898 60826 507134
rect 61062 506898 61146 507134
rect 61382 506898 61414 507134
rect 60794 471454 61414 506898
rect 60794 471218 60826 471454
rect 61062 471218 61146 471454
rect 61382 471218 61414 471454
rect 60794 471134 61414 471218
rect 60794 470898 60826 471134
rect 61062 470898 61146 471134
rect 61382 470898 61414 471134
rect 60794 435454 61414 470898
rect 60794 435218 60826 435454
rect 61062 435218 61146 435454
rect 61382 435218 61414 435454
rect 60794 435134 61414 435218
rect 60794 434898 60826 435134
rect 61062 434898 61146 435134
rect 61382 434898 61414 435134
rect 60794 399454 61414 434898
rect 60794 399218 60826 399454
rect 61062 399218 61146 399454
rect 61382 399218 61414 399454
rect 60794 399134 61414 399218
rect 60794 398898 60826 399134
rect 61062 398898 61146 399134
rect 61382 398898 61414 399134
rect 60794 363454 61414 398898
rect 60794 363218 60826 363454
rect 61062 363218 61146 363454
rect 61382 363218 61414 363454
rect 60794 363134 61414 363218
rect 60794 362898 60826 363134
rect 61062 362898 61146 363134
rect 61382 362898 61414 363134
rect 60794 327454 61414 362898
rect 60794 327218 60826 327454
rect 61062 327218 61146 327454
rect 61382 327218 61414 327454
rect 60794 327134 61414 327218
rect 60794 326898 60826 327134
rect 61062 326898 61146 327134
rect 61382 326898 61414 327134
rect 60794 291454 61414 326898
rect 60794 291218 60826 291454
rect 61062 291218 61146 291454
rect 61382 291218 61414 291454
rect 60794 291134 61414 291218
rect 60794 290898 60826 291134
rect 61062 290898 61146 291134
rect 61382 290898 61414 291134
rect 60794 255454 61414 290898
rect 60794 255218 60826 255454
rect 61062 255218 61146 255454
rect 61382 255218 61414 255454
rect 60794 255134 61414 255218
rect 60794 254898 60826 255134
rect 61062 254898 61146 255134
rect 61382 254898 61414 255134
rect 60794 219454 61414 254898
rect 60794 219218 60826 219454
rect 61062 219218 61146 219454
rect 61382 219218 61414 219454
rect 60794 219134 61414 219218
rect 60794 218898 60826 219134
rect 61062 218898 61146 219134
rect 61382 218898 61414 219134
rect 60794 183454 61414 218898
rect 60794 183218 60826 183454
rect 61062 183218 61146 183454
rect 61382 183218 61414 183454
rect 60794 183134 61414 183218
rect 60794 182898 60826 183134
rect 61062 182898 61146 183134
rect 61382 182898 61414 183134
rect 60794 147454 61414 182898
rect 60794 147218 60826 147454
rect 61062 147218 61146 147454
rect 61382 147218 61414 147454
rect 60794 147134 61414 147218
rect 60794 146898 60826 147134
rect 61062 146898 61146 147134
rect 61382 146898 61414 147134
rect 60794 111454 61414 146898
rect 60794 111218 60826 111454
rect 61062 111218 61146 111454
rect 61382 111218 61414 111454
rect 60794 111134 61414 111218
rect 60794 110898 60826 111134
rect 61062 110898 61146 111134
rect 61382 110898 61414 111134
rect 60794 75454 61414 110898
rect 60794 75218 60826 75454
rect 61062 75218 61146 75454
rect 61382 75218 61414 75454
rect 60794 75134 61414 75218
rect 60794 74898 60826 75134
rect 61062 74898 61146 75134
rect 61382 74898 61414 75134
rect 60794 74295 61414 74898
rect 61954 680614 62574 711002
rect 71954 710598 72574 711590
rect 71954 710362 71986 710598
rect 72222 710362 72306 710598
rect 72542 710362 72574 710598
rect 71954 710278 72574 710362
rect 71954 710042 71986 710278
rect 72222 710042 72306 710278
rect 72542 710042 72574 710278
rect 68234 708678 68854 709670
rect 68234 708442 68266 708678
rect 68502 708442 68586 708678
rect 68822 708442 68854 708678
rect 68234 708358 68854 708442
rect 68234 708122 68266 708358
rect 68502 708122 68586 708358
rect 68822 708122 68854 708358
rect 61954 680378 61986 680614
rect 62222 680378 62306 680614
rect 62542 680378 62574 680614
rect 61954 680294 62574 680378
rect 61954 680058 61986 680294
rect 62222 680058 62306 680294
rect 62542 680058 62574 680294
rect 61954 644614 62574 680058
rect 61954 644378 61986 644614
rect 62222 644378 62306 644614
rect 62542 644378 62574 644614
rect 61954 644294 62574 644378
rect 61954 644058 61986 644294
rect 62222 644058 62306 644294
rect 62542 644058 62574 644294
rect 61954 608614 62574 644058
rect 61954 608378 61986 608614
rect 62222 608378 62306 608614
rect 62542 608378 62574 608614
rect 61954 608294 62574 608378
rect 61954 608058 61986 608294
rect 62222 608058 62306 608294
rect 62542 608058 62574 608294
rect 61954 572614 62574 608058
rect 61954 572378 61986 572614
rect 62222 572378 62306 572614
rect 62542 572378 62574 572614
rect 61954 572294 62574 572378
rect 61954 572058 61986 572294
rect 62222 572058 62306 572294
rect 62542 572058 62574 572294
rect 61954 536614 62574 572058
rect 61954 536378 61986 536614
rect 62222 536378 62306 536614
rect 62542 536378 62574 536614
rect 61954 536294 62574 536378
rect 61954 536058 61986 536294
rect 62222 536058 62306 536294
rect 62542 536058 62574 536294
rect 61954 500614 62574 536058
rect 61954 500378 61986 500614
rect 62222 500378 62306 500614
rect 62542 500378 62574 500614
rect 61954 500294 62574 500378
rect 61954 500058 61986 500294
rect 62222 500058 62306 500294
rect 62542 500058 62574 500294
rect 61954 464614 62574 500058
rect 61954 464378 61986 464614
rect 62222 464378 62306 464614
rect 62542 464378 62574 464614
rect 61954 464294 62574 464378
rect 61954 464058 61986 464294
rect 62222 464058 62306 464294
rect 62542 464058 62574 464294
rect 61954 428614 62574 464058
rect 61954 428378 61986 428614
rect 62222 428378 62306 428614
rect 62542 428378 62574 428614
rect 61954 428294 62574 428378
rect 61954 428058 61986 428294
rect 62222 428058 62306 428294
rect 62542 428058 62574 428294
rect 61954 392614 62574 428058
rect 61954 392378 61986 392614
rect 62222 392378 62306 392614
rect 62542 392378 62574 392614
rect 61954 392294 62574 392378
rect 61954 392058 61986 392294
rect 62222 392058 62306 392294
rect 62542 392058 62574 392294
rect 61954 356614 62574 392058
rect 61954 356378 61986 356614
rect 62222 356378 62306 356614
rect 62542 356378 62574 356614
rect 61954 356294 62574 356378
rect 61954 356058 61986 356294
rect 62222 356058 62306 356294
rect 62542 356058 62574 356294
rect 61954 320614 62574 356058
rect 61954 320378 61986 320614
rect 62222 320378 62306 320614
rect 62542 320378 62574 320614
rect 61954 320294 62574 320378
rect 61954 320058 61986 320294
rect 62222 320058 62306 320294
rect 62542 320058 62574 320294
rect 61954 284614 62574 320058
rect 61954 284378 61986 284614
rect 62222 284378 62306 284614
rect 62542 284378 62574 284614
rect 61954 284294 62574 284378
rect 61954 284058 61986 284294
rect 62222 284058 62306 284294
rect 62542 284058 62574 284294
rect 61954 248614 62574 284058
rect 61954 248378 61986 248614
rect 62222 248378 62306 248614
rect 62542 248378 62574 248614
rect 61954 248294 62574 248378
rect 61954 248058 61986 248294
rect 62222 248058 62306 248294
rect 62542 248058 62574 248294
rect 61954 212614 62574 248058
rect 61954 212378 61986 212614
rect 62222 212378 62306 212614
rect 62542 212378 62574 212614
rect 61954 212294 62574 212378
rect 61954 212058 61986 212294
rect 62222 212058 62306 212294
rect 62542 212058 62574 212294
rect 61954 176614 62574 212058
rect 61954 176378 61986 176614
rect 62222 176378 62306 176614
rect 62542 176378 62574 176614
rect 61954 176294 62574 176378
rect 61954 176058 61986 176294
rect 62222 176058 62306 176294
rect 62542 176058 62574 176294
rect 61954 140614 62574 176058
rect 61954 140378 61986 140614
rect 62222 140378 62306 140614
rect 62542 140378 62574 140614
rect 61954 140294 62574 140378
rect 61954 140058 61986 140294
rect 62222 140058 62306 140294
rect 62542 140058 62574 140294
rect 61954 104614 62574 140058
rect 61954 104378 61986 104614
rect 62222 104378 62306 104614
rect 62542 104378 62574 104614
rect 61954 104294 62574 104378
rect 61954 104058 61986 104294
rect 62222 104058 62306 104294
rect 62542 104058 62574 104294
rect 61954 74295 62574 104058
rect 64514 706758 65134 707750
rect 64514 706522 64546 706758
rect 64782 706522 64866 706758
rect 65102 706522 65134 706758
rect 64514 706438 65134 706522
rect 64514 706202 64546 706438
rect 64782 706202 64866 706438
rect 65102 706202 65134 706438
rect 64514 691174 65134 706202
rect 64514 690938 64546 691174
rect 64782 690938 64866 691174
rect 65102 690938 65134 691174
rect 64514 690854 65134 690938
rect 64514 690618 64546 690854
rect 64782 690618 64866 690854
rect 65102 690618 65134 690854
rect 64514 655174 65134 690618
rect 64514 654938 64546 655174
rect 64782 654938 64866 655174
rect 65102 654938 65134 655174
rect 64514 654854 65134 654938
rect 64514 654618 64546 654854
rect 64782 654618 64866 654854
rect 65102 654618 65134 654854
rect 64514 619174 65134 654618
rect 64514 618938 64546 619174
rect 64782 618938 64866 619174
rect 65102 618938 65134 619174
rect 64514 618854 65134 618938
rect 64514 618618 64546 618854
rect 64782 618618 64866 618854
rect 65102 618618 65134 618854
rect 64514 583174 65134 618618
rect 64514 582938 64546 583174
rect 64782 582938 64866 583174
rect 65102 582938 65134 583174
rect 64514 582854 65134 582938
rect 64514 582618 64546 582854
rect 64782 582618 64866 582854
rect 65102 582618 65134 582854
rect 64514 547174 65134 582618
rect 64514 546938 64546 547174
rect 64782 546938 64866 547174
rect 65102 546938 65134 547174
rect 64514 546854 65134 546938
rect 64514 546618 64546 546854
rect 64782 546618 64866 546854
rect 65102 546618 65134 546854
rect 64514 511174 65134 546618
rect 64514 510938 64546 511174
rect 64782 510938 64866 511174
rect 65102 510938 65134 511174
rect 64514 510854 65134 510938
rect 64514 510618 64546 510854
rect 64782 510618 64866 510854
rect 65102 510618 65134 510854
rect 64514 475174 65134 510618
rect 64514 474938 64546 475174
rect 64782 474938 64866 475174
rect 65102 474938 65134 475174
rect 64514 474854 65134 474938
rect 64514 474618 64546 474854
rect 64782 474618 64866 474854
rect 65102 474618 65134 474854
rect 64514 439174 65134 474618
rect 64514 438938 64546 439174
rect 64782 438938 64866 439174
rect 65102 438938 65134 439174
rect 64514 438854 65134 438938
rect 64514 438618 64546 438854
rect 64782 438618 64866 438854
rect 65102 438618 65134 438854
rect 64514 403174 65134 438618
rect 64514 402938 64546 403174
rect 64782 402938 64866 403174
rect 65102 402938 65134 403174
rect 64514 402854 65134 402938
rect 64514 402618 64546 402854
rect 64782 402618 64866 402854
rect 65102 402618 65134 402854
rect 64514 367174 65134 402618
rect 64514 366938 64546 367174
rect 64782 366938 64866 367174
rect 65102 366938 65134 367174
rect 64514 366854 65134 366938
rect 64514 366618 64546 366854
rect 64782 366618 64866 366854
rect 65102 366618 65134 366854
rect 64514 331174 65134 366618
rect 64514 330938 64546 331174
rect 64782 330938 64866 331174
rect 65102 330938 65134 331174
rect 64514 330854 65134 330938
rect 64514 330618 64546 330854
rect 64782 330618 64866 330854
rect 65102 330618 65134 330854
rect 64514 295174 65134 330618
rect 64514 294938 64546 295174
rect 64782 294938 64866 295174
rect 65102 294938 65134 295174
rect 64514 294854 65134 294938
rect 64514 294618 64546 294854
rect 64782 294618 64866 294854
rect 65102 294618 65134 294854
rect 64514 259174 65134 294618
rect 64514 258938 64546 259174
rect 64782 258938 64866 259174
rect 65102 258938 65134 259174
rect 64514 258854 65134 258938
rect 64514 258618 64546 258854
rect 64782 258618 64866 258854
rect 65102 258618 65134 258854
rect 64514 223174 65134 258618
rect 64514 222938 64546 223174
rect 64782 222938 64866 223174
rect 65102 222938 65134 223174
rect 64514 222854 65134 222938
rect 64514 222618 64546 222854
rect 64782 222618 64866 222854
rect 65102 222618 65134 222854
rect 64514 187174 65134 222618
rect 64514 186938 64546 187174
rect 64782 186938 64866 187174
rect 65102 186938 65134 187174
rect 64514 186854 65134 186938
rect 64514 186618 64546 186854
rect 64782 186618 64866 186854
rect 65102 186618 65134 186854
rect 64514 151174 65134 186618
rect 64514 150938 64546 151174
rect 64782 150938 64866 151174
rect 65102 150938 65134 151174
rect 64514 150854 65134 150938
rect 64514 150618 64546 150854
rect 64782 150618 64866 150854
rect 65102 150618 65134 150854
rect 64514 115174 65134 150618
rect 64514 114938 64546 115174
rect 64782 114938 64866 115174
rect 65102 114938 65134 115174
rect 64514 114854 65134 114938
rect 64514 114618 64546 114854
rect 64782 114618 64866 114854
rect 65102 114618 65134 114854
rect 64514 79174 65134 114618
rect 64514 78938 64546 79174
rect 64782 78938 64866 79174
rect 65102 78938 65134 79174
rect 64514 78854 65134 78938
rect 64514 78618 64546 78854
rect 64782 78618 64866 78854
rect 65102 78618 65134 78854
rect 64514 74295 65134 78618
rect 68234 694894 68854 708122
rect 68234 694658 68266 694894
rect 68502 694658 68586 694894
rect 68822 694658 68854 694894
rect 68234 694574 68854 694658
rect 68234 694338 68266 694574
rect 68502 694338 68586 694574
rect 68822 694338 68854 694574
rect 68234 658894 68854 694338
rect 68234 658658 68266 658894
rect 68502 658658 68586 658894
rect 68822 658658 68854 658894
rect 68234 658574 68854 658658
rect 68234 658338 68266 658574
rect 68502 658338 68586 658574
rect 68822 658338 68854 658574
rect 68234 622894 68854 658338
rect 68234 622658 68266 622894
rect 68502 622658 68586 622894
rect 68822 622658 68854 622894
rect 68234 622574 68854 622658
rect 68234 622338 68266 622574
rect 68502 622338 68586 622574
rect 68822 622338 68854 622574
rect 68234 586894 68854 622338
rect 68234 586658 68266 586894
rect 68502 586658 68586 586894
rect 68822 586658 68854 586894
rect 68234 586574 68854 586658
rect 68234 586338 68266 586574
rect 68502 586338 68586 586574
rect 68822 586338 68854 586574
rect 68234 550894 68854 586338
rect 68234 550658 68266 550894
rect 68502 550658 68586 550894
rect 68822 550658 68854 550894
rect 68234 550574 68854 550658
rect 68234 550338 68266 550574
rect 68502 550338 68586 550574
rect 68822 550338 68854 550574
rect 68234 514894 68854 550338
rect 68234 514658 68266 514894
rect 68502 514658 68586 514894
rect 68822 514658 68854 514894
rect 68234 514574 68854 514658
rect 68234 514338 68266 514574
rect 68502 514338 68586 514574
rect 68822 514338 68854 514574
rect 68234 478894 68854 514338
rect 68234 478658 68266 478894
rect 68502 478658 68586 478894
rect 68822 478658 68854 478894
rect 68234 478574 68854 478658
rect 68234 478338 68266 478574
rect 68502 478338 68586 478574
rect 68822 478338 68854 478574
rect 68234 442894 68854 478338
rect 68234 442658 68266 442894
rect 68502 442658 68586 442894
rect 68822 442658 68854 442894
rect 68234 442574 68854 442658
rect 68234 442338 68266 442574
rect 68502 442338 68586 442574
rect 68822 442338 68854 442574
rect 68234 406894 68854 442338
rect 68234 406658 68266 406894
rect 68502 406658 68586 406894
rect 68822 406658 68854 406894
rect 68234 406574 68854 406658
rect 68234 406338 68266 406574
rect 68502 406338 68586 406574
rect 68822 406338 68854 406574
rect 68234 370894 68854 406338
rect 68234 370658 68266 370894
rect 68502 370658 68586 370894
rect 68822 370658 68854 370894
rect 68234 370574 68854 370658
rect 68234 370338 68266 370574
rect 68502 370338 68586 370574
rect 68822 370338 68854 370574
rect 68234 334894 68854 370338
rect 68234 334658 68266 334894
rect 68502 334658 68586 334894
rect 68822 334658 68854 334894
rect 68234 334574 68854 334658
rect 68234 334338 68266 334574
rect 68502 334338 68586 334574
rect 68822 334338 68854 334574
rect 68234 298894 68854 334338
rect 68234 298658 68266 298894
rect 68502 298658 68586 298894
rect 68822 298658 68854 298894
rect 68234 298574 68854 298658
rect 68234 298338 68266 298574
rect 68502 298338 68586 298574
rect 68822 298338 68854 298574
rect 68234 262894 68854 298338
rect 68234 262658 68266 262894
rect 68502 262658 68586 262894
rect 68822 262658 68854 262894
rect 68234 262574 68854 262658
rect 68234 262338 68266 262574
rect 68502 262338 68586 262574
rect 68822 262338 68854 262574
rect 68234 226894 68854 262338
rect 68234 226658 68266 226894
rect 68502 226658 68586 226894
rect 68822 226658 68854 226894
rect 68234 226574 68854 226658
rect 68234 226338 68266 226574
rect 68502 226338 68586 226574
rect 68822 226338 68854 226574
rect 68234 190894 68854 226338
rect 68234 190658 68266 190894
rect 68502 190658 68586 190894
rect 68822 190658 68854 190894
rect 68234 190574 68854 190658
rect 68234 190338 68266 190574
rect 68502 190338 68586 190574
rect 68822 190338 68854 190574
rect 68234 154894 68854 190338
rect 68234 154658 68266 154894
rect 68502 154658 68586 154894
rect 68822 154658 68854 154894
rect 68234 154574 68854 154658
rect 68234 154338 68266 154574
rect 68502 154338 68586 154574
rect 68822 154338 68854 154574
rect 68234 118894 68854 154338
rect 68234 118658 68266 118894
rect 68502 118658 68586 118894
rect 68822 118658 68854 118894
rect 68234 118574 68854 118658
rect 68234 118338 68266 118574
rect 68502 118338 68586 118574
rect 68822 118338 68854 118574
rect 68234 82894 68854 118338
rect 68234 82658 68266 82894
rect 68502 82658 68586 82894
rect 68822 82658 68854 82894
rect 68234 82574 68854 82658
rect 68234 82338 68266 82574
rect 68502 82338 68586 82574
rect 68822 82338 68854 82574
rect 68234 74295 68854 82338
rect 70794 705798 71414 705830
rect 70794 705562 70826 705798
rect 71062 705562 71146 705798
rect 71382 705562 71414 705798
rect 70794 705478 71414 705562
rect 70794 705242 70826 705478
rect 71062 705242 71146 705478
rect 71382 705242 71414 705478
rect 70794 669454 71414 705242
rect 70794 669218 70826 669454
rect 71062 669218 71146 669454
rect 71382 669218 71414 669454
rect 70794 669134 71414 669218
rect 70794 668898 70826 669134
rect 71062 668898 71146 669134
rect 71382 668898 71414 669134
rect 70794 633454 71414 668898
rect 70794 633218 70826 633454
rect 71062 633218 71146 633454
rect 71382 633218 71414 633454
rect 70794 633134 71414 633218
rect 70794 632898 70826 633134
rect 71062 632898 71146 633134
rect 71382 632898 71414 633134
rect 70794 597454 71414 632898
rect 70794 597218 70826 597454
rect 71062 597218 71146 597454
rect 71382 597218 71414 597454
rect 70794 597134 71414 597218
rect 70794 596898 70826 597134
rect 71062 596898 71146 597134
rect 71382 596898 71414 597134
rect 70794 561454 71414 596898
rect 70794 561218 70826 561454
rect 71062 561218 71146 561454
rect 71382 561218 71414 561454
rect 70794 561134 71414 561218
rect 70794 560898 70826 561134
rect 71062 560898 71146 561134
rect 71382 560898 71414 561134
rect 70794 525454 71414 560898
rect 70794 525218 70826 525454
rect 71062 525218 71146 525454
rect 71382 525218 71414 525454
rect 70794 525134 71414 525218
rect 70794 524898 70826 525134
rect 71062 524898 71146 525134
rect 71382 524898 71414 525134
rect 70794 489454 71414 524898
rect 70794 489218 70826 489454
rect 71062 489218 71146 489454
rect 71382 489218 71414 489454
rect 70794 489134 71414 489218
rect 70794 488898 70826 489134
rect 71062 488898 71146 489134
rect 71382 488898 71414 489134
rect 70794 453454 71414 488898
rect 70794 453218 70826 453454
rect 71062 453218 71146 453454
rect 71382 453218 71414 453454
rect 70794 453134 71414 453218
rect 70794 452898 70826 453134
rect 71062 452898 71146 453134
rect 71382 452898 71414 453134
rect 70794 417454 71414 452898
rect 70794 417218 70826 417454
rect 71062 417218 71146 417454
rect 71382 417218 71414 417454
rect 70794 417134 71414 417218
rect 70794 416898 70826 417134
rect 71062 416898 71146 417134
rect 71382 416898 71414 417134
rect 70794 381454 71414 416898
rect 70794 381218 70826 381454
rect 71062 381218 71146 381454
rect 71382 381218 71414 381454
rect 70794 381134 71414 381218
rect 70794 380898 70826 381134
rect 71062 380898 71146 381134
rect 71382 380898 71414 381134
rect 70794 345454 71414 380898
rect 70794 345218 70826 345454
rect 71062 345218 71146 345454
rect 71382 345218 71414 345454
rect 70794 345134 71414 345218
rect 70794 344898 70826 345134
rect 71062 344898 71146 345134
rect 71382 344898 71414 345134
rect 70794 309454 71414 344898
rect 70794 309218 70826 309454
rect 71062 309218 71146 309454
rect 71382 309218 71414 309454
rect 70794 309134 71414 309218
rect 70794 308898 70826 309134
rect 71062 308898 71146 309134
rect 71382 308898 71414 309134
rect 70794 273454 71414 308898
rect 70794 273218 70826 273454
rect 71062 273218 71146 273454
rect 71382 273218 71414 273454
rect 70794 273134 71414 273218
rect 70794 272898 70826 273134
rect 71062 272898 71146 273134
rect 71382 272898 71414 273134
rect 70794 237454 71414 272898
rect 70794 237218 70826 237454
rect 71062 237218 71146 237454
rect 71382 237218 71414 237454
rect 70794 237134 71414 237218
rect 70794 236898 70826 237134
rect 71062 236898 71146 237134
rect 71382 236898 71414 237134
rect 70794 201454 71414 236898
rect 70794 201218 70826 201454
rect 71062 201218 71146 201454
rect 71382 201218 71414 201454
rect 70794 201134 71414 201218
rect 70794 200898 70826 201134
rect 71062 200898 71146 201134
rect 71382 200898 71414 201134
rect 70794 165454 71414 200898
rect 70794 165218 70826 165454
rect 71062 165218 71146 165454
rect 71382 165218 71414 165454
rect 70794 165134 71414 165218
rect 70794 164898 70826 165134
rect 71062 164898 71146 165134
rect 71382 164898 71414 165134
rect 70794 129454 71414 164898
rect 70794 129218 70826 129454
rect 71062 129218 71146 129454
rect 71382 129218 71414 129454
rect 70794 129134 71414 129218
rect 70794 128898 70826 129134
rect 71062 128898 71146 129134
rect 71382 128898 71414 129134
rect 70794 93454 71414 128898
rect 70794 93218 70826 93454
rect 71062 93218 71146 93454
rect 71382 93218 71414 93454
rect 70794 93134 71414 93218
rect 70794 92898 70826 93134
rect 71062 92898 71146 93134
rect 71382 92898 71414 93134
rect 70794 74295 71414 92898
rect 71954 698614 72574 710042
rect 81954 711558 82574 711590
rect 81954 711322 81986 711558
rect 82222 711322 82306 711558
rect 82542 711322 82574 711558
rect 81954 711238 82574 711322
rect 81954 711002 81986 711238
rect 82222 711002 82306 711238
rect 82542 711002 82574 711238
rect 78234 709638 78854 709670
rect 78234 709402 78266 709638
rect 78502 709402 78586 709638
rect 78822 709402 78854 709638
rect 78234 709318 78854 709402
rect 78234 709082 78266 709318
rect 78502 709082 78586 709318
rect 78822 709082 78854 709318
rect 71954 698378 71986 698614
rect 72222 698378 72306 698614
rect 72542 698378 72574 698614
rect 71954 698294 72574 698378
rect 71954 698058 71986 698294
rect 72222 698058 72306 698294
rect 72542 698058 72574 698294
rect 71954 662614 72574 698058
rect 71954 662378 71986 662614
rect 72222 662378 72306 662614
rect 72542 662378 72574 662614
rect 71954 662294 72574 662378
rect 71954 662058 71986 662294
rect 72222 662058 72306 662294
rect 72542 662058 72574 662294
rect 71954 626614 72574 662058
rect 71954 626378 71986 626614
rect 72222 626378 72306 626614
rect 72542 626378 72574 626614
rect 71954 626294 72574 626378
rect 71954 626058 71986 626294
rect 72222 626058 72306 626294
rect 72542 626058 72574 626294
rect 71954 590614 72574 626058
rect 71954 590378 71986 590614
rect 72222 590378 72306 590614
rect 72542 590378 72574 590614
rect 71954 590294 72574 590378
rect 71954 590058 71986 590294
rect 72222 590058 72306 590294
rect 72542 590058 72574 590294
rect 71954 554614 72574 590058
rect 71954 554378 71986 554614
rect 72222 554378 72306 554614
rect 72542 554378 72574 554614
rect 71954 554294 72574 554378
rect 71954 554058 71986 554294
rect 72222 554058 72306 554294
rect 72542 554058 72574 554294
rect 71954 518614 72574 554058
rect 71954 518378 71986 518614
rect 72222 518378 72306 518614
rect 72542 518378 72574 518614
rect 71954 518294 72574 518378
rect 71954 518058 71986 518294
rect 72222 518058 72306 518294
rect 72542 518058 72574 518294
rect 71954 482614 72574 518058
rect 71954 482378 71986 482614
rect 72222 482378 72306 482614
rect 72542 482378 72574 482614
rect 71954 482294 72574 482378
rect 71954 482058 71986 482294
rect 72222 482058 72306 482294
rect 72542 482058 72574 482294
rect 71954 446614 72574 482058
rect 71954 446378 71986 446614
rect 72222 446378 72306 446614
rect 72542 446378 72574 446614
rect 71954 446294 72574 446378
rect 71954 446058 71986 446294
rect 72222 446058 72306 446294
rect 72542 446058 72574 446294
rect 71954 410614 72574 446058
rect 71954 410378 71986 410614
rect 72222 410378 72306 410614
rect 72542 410378 72574 410614
rect 71954 410294 72574 410378
rect 71954 410058 71986 410294
rect 72222 410058 72306 410294
rect 72542 410058 72574 410294
rect 71954 374614 72574 410058
rect 71954 374378 71986 374614
rect 72222 374378 72306 374614
rect 72542 374378 72574 374614
rect 71954 374294 72574 374378
rect 71954 374058 71986 374294
rect 72222 374058 72306 374294
rect 72542 374058 72574 374294
rect 71954 338614 72574 374058
rect 71954 338378 71986 338614
rect 72222 338378 72306 338614
rect 72542 338378 72574 338614
rect 71954 338294 72574 338378
rect 71954 338058 71986 338294
rect 72222 338058 72306 338294
rect 72542 338058 72574 338294
rect 71954 302614 72574 338058
rect 71954 302378 71986 302614
rect 72222 302378 72306 302614
rect 72542 302378 72574 302614
rect 71954 302294 72574 302378
rect 71954 302058 71986 302294
rect 72222 302058 72306 302294
rect 72542 302058 72574 302294
rect 71954 266614 72574 302058
rect 71954 266378 71986 266614
rect 72222 266378 72306 266614
rect 72542 266378 72574 266614
rect 71954 266294 72574 266378
rect 71954 266058 71986 266294
rect 72222 266058 72306 266294
rect 72542 266058 72574 266294
rect 71954 230614 72574 266058
rect 71954 230378 71986 230614
rect 72222 230378 72306 230614
rect 72542 230378 72574 230614
rect 71954 230294 72574 230378
rect 71954 230058 71986 230294
rect 72222 230058 72306 230294
rect 72542 230058 72574 230294
rect 71954 194614 72574 230058
rect 71954 194378 71986 194614
rect 72222 194378 72306 194614
rect 72542 194378 72574 194614
rect 71954 194294 72574 194378
rect 71954 194058 71986 194294
rect 72222 194058 72306 194294
rect 72542 194058 72574 194294
rect 71954 158614 72574 194058
rect 71954 158378 71986 158614
rect 72222 158378 72306 158614
rect 72542 158378 72574 158614
rect 71954 158294 72574 158378
rect 71954 158058 71986 158294
rect 72222 158058 72306 158294
rect 72542 158058 72574 158294
rect 71954 122614 72574 158058
rect 71954 122378 71986 122614
rect 72222 122378 72306 122614
rect 72542 122378 72574 122614
rect 71954 122294 72574 122378
rect 71954 122058 71986 122294
rect 72222 122058 72306 122294
rect 72542 122058 72574 122294
rect 71954 86614 72574 122058
rect 71954 86378 71986 86614
rect 72222 86378 72306 86614
rect 72542 86378 72574 86614
rect 71954 86294 72574 86378
rect 71954 86058 71986 86294
rect 72222 86058 72306 86294
rect 72542 86058 72574 86294
rect 71954 74295 72574 86058
rect 74514 707718 75134 707750
rect 74514 707482 74546 707718
rect 74782 707482 74866 707718
rect 75102 707482 75134 707718
rect 74514 707398 75134 707482
rect 74514 707162 74546 707398
rect 74782 707162 74866 707398
rect 75102 707162 75134 707398
rect 74514 673174 75134 707162
rect 74514 672938 74546 673174
rect 74782 672938 74866 673174
rect 75102 672938 75134 673174
rect 74514 672854 75134 672938
rect 74514 672618 74546 672854
rect 74782 672618 74866 672854
rect 75102 672618 75134 672854
rect 74514 637174 75134 672618
rect 74514 636938 74546 637174
rect 74782 636938 74866 637174
rect 75102 636938 75134 637174
rect 74514 636854 75134 636938
rect 74514 636618 74546 636854
rect 74782 636618 74866 636854
rect 75102 636618 75134 636854
rect 74514 601174 75134 636618
rect 74514 600938 74546 601174
rect 74782 600938 74866 601174
rect 75102 600938 75134 601174
rect 74514 600854 75134 600938
rect 74514 600618 74546 600854
rect 74782 600618 74866 600854
rect 75102 600618 75134 600854
rect 74514 565174 75134 600618
rect 74514 564938 74546 565174
rect 74782 564938 74866 565174
rect 75102 564938 75134 565174
rect 74514 564854 75134 564938
rect 74514 564618 74546 564854
rect 74782 564618 74866 564854
rect 75102 564618 75134 564854
rect 74514 529174 75134 564618
rect 74514 528938 74546 529174
rect 74782 528938 74866 529174
rect 75102 528938 75134 529174
rect 74514 528854 75134 528938
rect 74514 528618 74546 528854
rect 74782 528618 74866 528854
rect 75102 528618 75134 528854
rect 74514 493174 75134 528618
rect 74514 492938 74546 493174
rect 74782 492938 74866 493174
rect 75102 492938 75134 493174
rect 74514 492854 75134 492938
rect 74514 492618 74546 492854
rect 74782 492618 74866 492854
rect 75102 492618 75134 492854
rect 74514 457174 75134 492618
rect 74514 456938 74546 457174
rect 74782 456938 74866 457174
rect 75102 456938 75134 457174
rect 74514 456854 75134 456938
rect 74514 456618 74546 456854
rect 74782 456618 74866 456854
rect 75102 456618 75134 456854
rect 74514 421174 75134 456618
rect 74514 420938 74546 421174
rect 74782 420938 74866 421174
rect 75102 420938 75134 421174
rect 74514 420854 75134 420938
rect 74514 420618 74546 420854
rect 74782 420618 74866 420854
rect 75102 420618 75134 420854
rect 74514 385174 75134 420618
rect 74514 384938 74546 385174
rect 74782 384938 74866 385174
rect 75102 384938 75134 385174
rect 74514 384854 75134 384938
rect 74514 384618 74546 384854
rect 74782 384618 74866 384854
rect 75102 384618 75134 384854
rect 74514 349174 75134 384618
rect 74514 348938 74546 349174
rect 74782 348938 74866 349174
rect 75102 348938 75134 349174
rect 74514 348854 75134 348938
rect 74514 348618 74546 348854
rect 74782 348618 74866 348854
rect 75102 348618 75134 348854
rect 74514 313174 75134 348618
rect 74514 312938 74546 313174
rect 74782 312938 74866 313174
rect 75102 312938 75134 313174
rect 74514 312854 75134 312938
rect 74514 312618 74546 312854
rect 74782 312618 74866 312854
rect 75102 312618 75134 312854
rect 74514 277174 75134 312618
rect 74514 276938 74546 277174
rect 74782 276938 74866 277174
rect 75102 276938 75134 277174
rect 74514 276854 75134 276938
rect 74514 276618 74546 276854
rect 74782 276618 74866 276854
rect 75102 276618 75134 276854
rect 74514 241174 75134 276618
rect 74514 240938 74546 241174
rect 74782 240938 74866 241174
rect 75102 240938 75134 241174
rect 74514 240854 75134 240938
rect 74514 240618 74546 240854
rect 74782 240618 74866 240854
rect 75102 240618 75134 240854
rect 74514 205174 75134 240618
rect 74514 204938 74546 205174
rect 74782 204938 74866 205174
rect 75102 204938 75134 205174
rect 74514 204854 75134 204938
rect 74514 204618 74546 204854
rect 74782 204618 74866 204854
rect 75102 204618 75134 204854
rect 74514 169174 75134 204618
rect 74514 168938 74546 169174
rect 74782 168938 74866 169174
rect 75102 168938 75134 169174
rect 74514 168854 75134 168938
rect 74514 168618 74546 168854
rect 74782 168618 74866 168854
rect 75102 168618 75134 168854
rect 74514 133174 75134 168618
rect 74514 132938 74546 133174
rect 74782 132938 74866 133174
rect 75102 132938 75134 133174
rect 74514 132854 75134 132938
rect 74514 132618 74546 132854
rect 74782 132618 74866 132854
rect 75102 132618 75134 132854
rect 74514 97174 75134 132618
rect 74514 96938 74546 97174
rect 74782 96938 74866 97174
rect 75102 96938 75134 97174
rect 74514 96854 75134 96938
rect 74514 96618 74546 96854
rect 74782 96618 74866 96854
rect 75102 96618 75134 96854
rect 31523 71908 31589 71909
rect 31523 71844 31524 71908
rect 31588 71844 31589 71908
rect 31523 71843 31589 71844
rect 14514 60938 14546 61174
rect 14782 60938 14866 61174
rect 15102 60938 15134 61174
rect 14514 60854 15134 60938
rect 14514 60618 14546 60854
rect 14782 60618 14866 60854
rect 15102 60618 15134 60854
rect 14514 25174 15134 60618
rect 24208 39454 24528 39486
rect 24208 39218 24250 39454
rect 24486 39218 24528 39454
rect 24208 39134 24528 39218
rect 24208 38898 24250 39134
rect 24486 38898 24528 39134
rect 24208 38866 24528 38898
rect 14514 24938 14546 25174
rect 14782 24938 14866 25174
rect 15102 24938 15134 25174
rect 14514 24854 15134 24938
rect 14514 24618 14546 24854
rect 14782 24618 14866 24854
rect 15102 24618 15134 24854
rect 14514 -3226 15134 24618
rect 14514 -3462 14546 -3226
rect 14782 -3462 14866 -3226
rect 15102 -3462 15134 -3226
rect 14514 -3546 15134 -3462
rect 14514 -3782 14546 -3546
rect 14782 -3782 14866 -3546
rect 15102 -3782 15134 -3546
rect 14514 -3814 15134 -3782
rect 18234 -5146 18854 18000
rect 20794 3454 21414 18000
rect 20794 3218 20826 3454
rect 21062 3218 21146 3454
rect 21382 3218 21414 3454
rect 20794 3134 21414 3218
rect 20794 2898 20826 3134
rect 21062 2898 21146 3134
rect 21382 2898 21414 3134
rect 20794 -346 21414 2898
rect 20794 -582 20826 -346
rect 21062 -582 21146 -346
rect 21382 -582 21414 -346
rect 20794 -666 21414 -582
rect 20794 -902 20826 -666
rect 21062 -902 21146 -666
rect 21382 -902 21414 -666
rect 20794 -1894 21414 -902
rect 18234 -5382 18266 -5146
rect 18502 -5382 18586 -5146
rect 18822 -5382 18854 -5146
rect 18234 -5466 18854 -5382
rect 18234 -5702 18266 -5466
rect 18502 -5702 18586 -5466
rect 18822 -5702 18854 -5466
rect 18234 -5734 18854 -5702
rect 11954 -6342 11986 -6106
rect 12222 -6342 12306 -6106
rect 12542 -6342 12574 -6106
rect 11954 -6426 12574 -6342
rect 11954 -6662 11986 -6426
rect 12222 -6662 12306 -6426
rect 12542 -6662 12574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 11954 -7654 12574 -6662
rect 21954 -7066 22574 18000
rect 24514 7174 25134 18000
rect 24514 6938 24546 7174
rect 24782 6938 24866 7174
rect 25102 6938 25134 7174
rect 24514 6854 25134 6938
rect 24514 6618 24546 6854
rect 24782 6618 24866 6854
rect 25102 6618 25134 6854
rect 24514 -2266 25134 6618
rect 24514 -2502 24546 -2266
rect 24782 -2502 24866 -2266
rect 25102 -2502 25134 -2266
rect 24514 -2586 25134 -2502
rect 24514 -2822 24546 -2586
rect 24782 -2822 24866 -2586
rect 25102 -2822 25134 -2586
rect 24514 -3814 25134 -2822
rect 28234 10894 28854 18000
rect 28234 10658 28266 10894
rect 28502 10658 28586 10894
rect 28822 10658 28854 10894
rect 28234 10574 28854 10658
rect 28234 10338 28266 10574
rect 28502 10338 28586 10574
rect 28822 10338 28854 10574
rect 28234 -4186 28854 10338
rect 30794 -1306 31414 18000
rect 31526 5677 31586 71843
rect 74514 61174 75134 96618
rect 74514 60938 74546 61174
rect 74782 60938 74866 61174
rect 75102 60938 75134 61174
rect 74514 60854 75134 60938
rect 74514 60618 74546 60854
rect 74782 60618 74866 60854
rect 75102 60618 75134 60854
rect 39568 57454 39888 57486
rect 39568 57218 39610 57454
rect 39846 57218 39888 57454
rect 39568 57134 39888 57218
rect 39568 56898 39610 57134
rect 39846 56898 39888 57134
rect 39568 56866 39888 56898
rect 54928 39454 55248 39486
rect 54928 39218 54970 39454
rect 55206 39218 55248 39454
rect 54928 39134 55248 39218
rect 54928 38898 54970 39134
rect 55206 38898 55248 39134
rect 54928 38866 55248 38898
rect 74514 25174 75134 60618
rect 74514 24938 74546 25174
rect 74782 24938 74866 25174
rect 75102 24938 75134 25174
rect 74514 24854 75134 24938
rect 74514 24618 74546 24854
rect 74782 24618 74866 24854
rect 75102 24618 75134 24854
rect 31954 14614 32574 18000
rect 31954 14378 31986 14614
rect 32222 14378 32306 14614
rect 32542 14378 32574 14614
rect 31954 14294 32574 14378
rect 31954 14058 31986 14294
rect 32222 14058 32306 14294
rect 32542 14058 32574 14294
rect 31523 5676 31589 5677
rect 31523 5612 31524 5676
rect 31588 5612 31589 5676
rect 31523 5611 31589 5612
rect 30794 -1542 30826 -1306
rect 31062 -1542 31146 -1306
rect 31382 -1542 31414 -1306
rect 30794 -1626 31414 -1542
rect 30794 -1862 30826 -1626
rect 31062 -1862 31146 -1626
rect 31382 -1862 31414 -1626
rect 30794 -1894 31414 -1862
rect 28234 -4422 28266 -4186
rect 28502 -4422 28586 -4186
rect 28822 -4422 28854 -4186
rect 28234 -4506 28854 -4422
rect 28234 -4742 28266 -4506
rect 28502 -4742 28586 -4506
rect 28822 -4742 28854 -4506
rect 28234 -5734 28854 -4742
rect 21954 -7302 21986 -7066
rect 22222 -7302 22306 -7066
rect 22542 -7302 22574 -7066
rect 21954 -7386 22574 -7302
rect 21954 -7622 21986 -7386
rect 22222 -7622 22306 -7386
rect 22542 -7622 22574 -7386
rect 21954 -7654 22574 -7622
rect 31954 -6106 32574 14058
rect 34514 -3226 35134 18000
rect 34514 -3462 34546 -3226
rect 34782 -3462 34866 -3226
rect 35102 -3462 35134 -3226
rect 34514 -3546 35134 -3462
rect 34514 -3782 34546 -3546
rect 34782 -3782 34866 -3546
rect 35102 -3782 35134 -3546
rect 34514 -3814 35134 -3782
rect 38234 -5146 38854 18000
rect 40794 3454 41414 18000
rect 40794 3218 40826 3454
rect 41062 3218 41146 3454
rect 41382 3218 41414 3454
rect 40794 3134 41414 3218
rect 40794 2898 40826 3134
rect 41062 2898 41146 3134
rect 41382 2898 41414 3134
rect 40794 -346 41414 2898
rect 40794 -582 40826 -346
rect 41062 -582 41146 -346
rect 41382 -582 41414 -346
rect 40794 -666 41414 -582
rect 40794 -902 40826 -666
rect 41062 -902 41146 -666
rect 41382 -902 41414 -666
rect 40794 -1894 41414 -902
rect 38234 -5382 38266 -5146
rect 38502 -5382 38586 -5146
rect 38822 -5382 38854 -5146
rect 38234 -5466 38854 -5382
rect 38234 -5702 38266 -5466
rect 38502 -5702 38586 -5466
rect 38822 -5702 38854 -5466
rect 38234 -5734 38854 -5702
rect 31954 -6342 31986 -6106
rect 32222 -6342 32306 -6106
rect 32542 -6342 32574 -6106
rect 31954 -6426 32574 -6342
rect 31954 -6662 31986 -6426
rect 32222 -6662 32306 -6426
rect 32542 -6662 32574 -6426
rect 31954 -7654 32574 -6662
rect 41954 -7066 42574 18000
rect 44514 7174 45134 18000
rect 44514 6938 44546 7174
rect 44782 6938 44866 7174
rect 45102 6938 45134 7174
rect 44514 6854 45134 6938
rect 44514 6618 44546 6854
rect 44782 6618 44866 6854
rect 45102 6618 45134 6854
rect 44514 -2266 45134 6618
rect 44514 -2502 44546 -2266
rect 44782 -2502 44866 -2266
rect 45102 -2502 45134 -2266
rect 44514 -2586 45134 -2502
rect 44514 -2822 44546 -2586
rect 44782 -2822 44866 -2586
rect 45102 -2822 45134 -2586
rect 44514 -3814 45134 -2822
rect 48234 10894 48854 18000
rect 48234 10658 48266 10894
rect 48502 10658 48586 10894
rect 48822 10658 48854 10894
rect 48234 10574 48854 10658
rect 48234 10338 48266 10574
rect 48502 10338 48586 10574
rect 48822 10338 48854 10574
rect 48234 -4186 48854 10338
rect 50794 -1306 51414 18000
rect 50794 -1542 50826 -1306
rect 51062 -1542 51146 -1306
rect 51382 -1542 51414 -1306
rect 50794 -1626 51414 -1542
rect 50794 -1862 50826 -1626
rect 51062 -1862 51146 -1626
rect 51382 -1862 51414 -1626
rect 50794 -1894 51414 -1862
rect 51954 14614 52574 18000
rect 51954 14378 51986 14614
rect 52222 14378 52306 14614
rect 52542 14378 52574 14614
rect 51954 14294 52574 14378
rect 51954 14058 51986 14294
rect 52222 14058 52306 14294
rect 52542 14058 52574 14294
rect 48234 -4422 48266 -4186
rect 48502 -4422 48586 -4186
rect 48822 -4422 48854 -4186
rect 48234 -4506 48854 -4422
rect 48234 -4742 48266 -4506
rect 48502 -4742 48586 -4506
rect 48822 -4742 48854 -4506
rect 48234 -5734 48854 -4742
rect 41954 -7302 41986 -7066
rect 42222 -7302 42306 -7066
rect 42542 -7302 42574 -7066
rect 41954 -7386 42574 -7302
rect 41954 -7622 41986 -7386
rect 42222 -7622 42306 -7386
rect 42542 -7622 42574 -7386
rect 41954 -7654 42574 -7622
rect 51954 -6106 52574 14058
rect 54514 -3226 55134 18000
rect 54514 -3462 54546 -3226
rect 54782 -3462 54866 -3226
rect 55102 -3462 55134 -3226
rect 54514 -3546 55134 -3462
rect 54514 -3782 54546 -3546
rect 54782 -3782 54866 -3546
rect 55102 -3782 55134 -3546
rect 54514 -3814 55134 -3782
rect 58234 -5146 58854 18000
rect 60794 3454 61414 18000
rect 60794 3218 60826 3454
rect 61062 3218 61146 3454
rect 61382 3218 61414 3454
rect 60794 3134 61414 3218
rect 60794 2898 60826 3134
rect 61062 2898 61146 3134
rect 61382 2898 61414 3134
rect 60794 -346 61414 2898
rect 60794 -582 60826 -346
rect 61062 -582 61146 -346
rect 61382 -582 61414 -346
rect 60794 -666 61414 -582
rect 60794 -902 60826 -666
rect 61062 -902 61146 -666
rect 61382 -902 61414 -666
rect 60794 -1894 61414 -902
rect 58234 -5382 58266 -5146
rect 58502 -5382 58586 -5146
rect 58822 -5382 58854 -5146
rect 58234 -5466 58854 -5382
rect 58234 -5702 58266 -5466
rect 58502 -5702 58586 -5466
rect 58822 -5702 58854 -5466
rect 58234 -5734 58854 -5702
rect 51954 -6342 51986 -6106
rect 52222 -6342 52306 -6106
rect 52542 -6342 52574 -6106
rect 51954 -6426 52574 -6342
rect 51954 -6662 51986 -6426
rect 52222 -6662 52306 -6426
rect 52542 -6662 52574 -6426
rect 51954 -7654 52574 -6662
rect 61954 -7066 62574 18000
rect 64514 7174 65134 18000
rect 64514 6938 64546 7174
rect 64782 6938 64866 7174
rect 65102 6938 65134 7174
rect 64514 6854 65134 6938
rect 64514 6618 64546 6854
rect 64782 6618 64866 6854
rect 65102 6618 65134 6854
rect 64514 -2266 65134 6618
rect 64514 -2502 64546 -2266
rect 64782 -2502 64866 -2266
rect 65102 -2502 65134 -2266
rect 64514 -2586 65134 -2502
rect 64514 -2822 64546 -2586
rect 64782 -2822 64866 -2586
rect 65102 -2822 65134 -2586
rect 64514 -3814 65134 -2822
rect 68234 10894 68854 18000
rect 68234 10658 68266 10894
rect 68502 10658 68586 10894
rect 68822 10658 68854 10894
rect 68234 10574 68854 10658
rect 68234 10338 68266 10574
rect 68502 10338 68586 10574
rect 68822 10338 68854 10574
rect 68234 -4186 68854 10338
rect 70794 -1306 71414 18000
rect 70794 -1542 70826 -1306
rect 71062 -1542 71146 -1306
rect 71382 -1542 71414 -1306
rect 70794 -1626 71414 -1542
rect 70794 -1862 70826 -1626
rect 71062 -1862 71146 -1626
rect 71382 -1862 71414 -1626
rect 70794 -1894 71414 -1862
rect 71954 14614 72574 18000
rect 71954 14378 71986 14614
rect 72222 14378 72306 14614
rect 72542 14378 72574 14614
rect 71954 14294 72574 14378
rect 71954 14058 71986 14294
rect 72222 14058 72306 14294
rect 72542 14058 72574 14294
rect 68234 -4422 68266 -4186
rect 68502 -4422 68586 -4186
rect 68822 -4422 68854 -4186
rect 68234 -4506 68854 -4422
rect 68234 -4742 68266 -4506
rect 68502 -4742 68586 -4506
rect 68822 -4742 68854 -4506
rect 68234 -5734 68854 -4742
rect 61954 -7302 61986 -7066
rect 62222 -7302 62306 -7066
rect 62542 -7302 62574 -7066
rect 61954 -7386 62574 -7302
rect 61954 -7622 61986 -7386
rect 62222 -7622 62306 -7386
rect 62542 -7622 62574 -7386
rect 61954 -7654 62574 -7622
rect 71954 -6106 72574 14058
rect 74514 -3226 75134 24618
rect 74514 -3462 74546 -3226
rect 74782 -3462 74866 -3226
rect 75102 -3462 75134 -3226
rect 74514 -3546 75134 -3462
rect 74514 -3782 74546 -3546
rect 74782 -3782 74866 -3546
rect 75102 -3782 75134 -3546
rect 74514 -3814 75134 -3782
rect 78234 676894 78854 709082
rect 78234 676658 78266 676894
rect 78502 676658 78586 676894
rect 78822 676658 78854 676894
rect 78234 676574 78854 676658
rect 78234 676338 78266 676574
rect 78502 676338 78586 676574
rect 78822 676338 78854 676574
rect 78234 640894 78854 676338
rect 78234 640658 78266 640894
rect 78502 640658 78586 640894
rect 78822 640658 78854 640894
rect 78234 640574 78854 640658
rect 78234 640338 78266 640574
rect 78502 640338 78586 640574
rect 78822 640338 78854 640574
rect 78234 604894 78854 640338
rect 78234 604658 78266 604894
rect 78502 604658 78586 604894
rect 78822 604658 78854 604894
rect 78234 604574 78854 604658
rect 78234 604338 78266 604574
rect 78502 604338 78586 604574
rect 78822 604338 78854 604574
rect 78234 568894 78854 604338
rect 78234 568658 78266 568894
rect 78502 568658 78586 568894
rect 78822 568658 78854 568894
rect 78234 568574 78854 568658
rect 78234 568338 78266 568574
rect 78502 568338 78586 568574
rect 78822 568338 78854 568574
rect 78234 532894 78854 568338
rect 78234 532658 78266 532894
rect 78502 532658 78586 532894
rect 78822 532658 78854 532894
rect 78234 532574 78854 532658
rect 78234 532338 78266 532574
rect 78502 532338 78586 532574
rect 78822 532338 78854 532574
rect 78234 496894 78854 532338
rect 78234 496658 78266 496894
rect 78502 496658 78586 496894
rect 78822 496658 78854 496894
rect 78234 496574 78854 496658
rect 78234 496338 78266 496574
rect 78502 496338 78586 496574
rect 78822 496338 78854 496574
rect 78234 460894 78854 496338
rect 78234 460658 78266 460894
rect 78502 460658 78586 460894
rect 78822 460658 78854 460894
rect 78234 460574 78854 460658
rect 78234 460338 78266 460574
rect 78502 460338 78586 460574
rect 78822 460338 78854 460574
rect 78234 424894 78854 460338
rect 78234 424658 78266 424894
rect 78502 424658 78586 424894
rect 78822 424658 78854 424894
rect 78234 424574 78854 424658
rect 78234 424338 78266 424574
rect 78502 424338 78586 424574
rect 78822 424338 78854 424574
rect 78234 388894 78854 424338
rect 78234 388658 78266 388894
rect 78502 388658 78586 388894
rect 78822 388658 78854 388894
rect 78234 388574 78854 388658
rect 78234 388338 78266 388574
rect 78502 388338 78586 388574
rect 78822 388338 78854 388574
rect 78234 352894 78854 388338
rect 78234 352658 78266 352894
rect 78502 352658 78586 352894
rect 78822 352658 78854 352894
rect 78234 352574 78854 352658
rect 78234 352338 78266 352574
rect 78502 352338 78586 352574
rect 78822 352338 78854 352574
rect 78234 316894 78854 352338
rect 78234 316658 78266 316894
rect 78502 316658 78586 316894
rect 78822 316658 78854 316894
rect 78234 316574 78854 316658
rect 78234 316338 78266 316574
rect 78502 316338 78586 316574
rect 78822 316338 78854 316574
rect 78234 280894 78854 316338
rect 78234 280658 78266 280894
rect 78502 280658 78586 280894
rect 78822 280658 78854 280894
rect 78234 280574 78854 280658
rect 78234 280338 78266 280574
rect 78502 280338 78586 280574
rect 78822 280338 78854 280574
rect 78234 244894 78854 280338
rect 78234 244658 78266 244894
rect 78502 244658 78586 244894
rect 78822 244658 78854 244894
rect 78234 244574 78854 244658
rect 78234 244338 78266 244574
rect 78502 244338 78586 244574
rect 78822 244338 78854 244574
rect 78234 208894 78854 244338
rect 78234 208658 78266 208894
rect 78502 208658 78586 208894
rect 78822 208658 78854 208894
rect 78234 208574 78854 208658
rect 78234 208338 78266 208574
rect 78502 208338 78586 208574
rect 78822 208338 78854 208574
rect 78234 172894 78854 208338
rect 78234 172658 78266 172894
rect 78502 172658 78586 172894
rect 78822 172658 78854 172894
rect 78234 172574 78854 172658
rect 78234 172338 78266 172574
rect 78502 172338 78586 172574
rect 78822 172338 78854 172574
rect 78234 136894 78854 172338
rect 78234 136658 78266 136894
rect 78502 136658 78586 136894
rect 78822 136658 78854 136894
rect 78234 136574 78854 136658
rect 78234 136338 78266 136574
rect 78502 136338 78586 136574
rect 78822 136338 78854 136574
rect 78234 100894 78854 136338
rect 78234 100658 78266 100894
rect 78502 100658 78586 100894
rect 78822 100658 78854 100894
rect 78234 100574 78854 100658
rect 78234 100338 78266 100574
rect 78502 100338 78586 100574
rect 78822 100338 78854 100574
rect 78234 64894 78854 100338
rect 78234 64658 78266 64894
rect 78502 64658 78586 64894
rect 78822 64658 78854 64894
rect 78234 64574 78854 64658
rect 78234 64338 78266 64574
rect 78502 64338 78586 64574
rect 78822 64338 78854 64574
rect 78234 28894 78854 64338
rect 78234 28658 78266 28894
rect 78502 28658 78586 28894
rect 78822 28658 78854 28894
rect 78234 28574 78854 28658
rect 78234 28338 78266 28574
rect 78502 28338 78586 28574
rect 78822 28338 78854 28574
rect 78234 -5146 78854 28338
rect 80794 704838 81414 705830
rect 80794 704602 80826 704838
rect 81062 704602 81146 704838
rect 81382 704602 81414 704838
rect 80794 704518 81414 704602
rect 80794 704282 80826 704518
rect 81062 704282 81146 704518
rect 81382 704282 81414 704518
rect 80794 687454 81414 704282
rect 80794 687218 80826 687454
rect 81062 687218 81146 687454
rect 81382 687218 81414 687454
rect 80794 687134 81414 687218
rect 80794 686898 80826 687134
rect 81062 686898 81146 687134
rect 81382 686898 81414 687134
rect 80794 651454 81414 686898
rect 80794 651218 80826 651454
rect 81062 651218 81146 651454
rect 81382 651218 81414 651454
rect 80794 651134 81414 651218
rect 80794 650898 80826 651134
rect 81062 650898 81146 651134
rect 81382 650898 81414 651134
rect 80794 615454 81414 650898
rect 80794 615218 80826 615454
rect 81062 615218 81146 615454
rect 81382 615218 81414 615454
rect 80794 615134 81414 615218
rect 80794 614898 80826 615134
rect 81062 614898 81146 615134
rect 81382 614898 81414 615134
rect 80794 579454 81414 614898
rect 80794 579218 80826 579454
rect 81062 579218 81146 579454
rect 81382 579218 81414 579454
rect 80794 579134 81414 579218
rect 80794 578898 80826 579134
rect 81062 578898 81146 579134
rect 81382 578898 81414 579134
rect 80794 543454 81414 578898
rect 80794 543218 80826 543454
rect 81062 543218 81146 543454
rect 81382 543218 81414 543454
rect 80794 543134 81414 543218
rect 80794 542898 80826 543134
rect 81062 542898 81146 543134
rect 81382 542898 81414 543134
rect 80794 507454 81414 542898
rect 80794 507218 80826 507454
rect 81062 507218 81146 507454
rect 81382 507218 81414 507454
rect 80794 507134 81414 507218
rect 80794 506898 80826 507134
rect 81062 506898 81146 507134
rect 81382 506898 81414 507134
rect 80794 471454 81414 506898
rect 80794 471218 80826 471454
rect 81062 471218 81146 471454
rect 81382 471218 81414 471454
rect 80794 471134 81414 471218
rect 80794 470898 80826 471134
rect 81062 470898 81146 471134
rect 81382 470898 81414 471134
rect 80794 435454 81414 470898
rect 80794 435218 80826 435454
rect 81062 435218 81146 435454
rect 81382 435218 81414 435454
rect 80794 435134 81414 435218
rect 80794 434898 80826 435134
rect 81062 434898 81146 435134
rect 81382 434898 81414 435134
rect 80794 399454 81414 434898
rect 80794 399218 80826 399454
rect 81062 399218 81146 399454
rect 81382 399218 81414 399454
rect 80794 399134 81414 399218
rect 80794 398898 80826 399134
rect 81062 398898 81146 399134
rect 81382 398898 81414 399134
rect 80794 363454 81414 398898
rect 80794 363218 80826 363454
rect 81062 363218 81146 363454
rect 81382 363218 81414 363454
rect 80794 363134 81414 363218
rect 80794 362898 80826 363134
rect 81062 362898 81146 363134
rect 81382 362898 81414 363134
rect 80794 327454 81414 362898
rect 80794 327218 80826 327454
rect 81062 327218 81146 327454
rect 81382 327218 81414 327454
rect 80794 327134 81414 327218
rect 80794 326898 80826 327134
rect 81062 326898 81146 327134
rect 81382 326898 81414 327134
rect 80794 291454 81414 326898
rect 80794 291218 80826 291454
rect 81062 291218 81146 291454
rect 81382 291218 81414 291454
rect 80794 291134 81414 291218
rect 80794 290898 80826 291134
rect 81062 290898 81146 291134
rect 81382 290898 81414 291134
rect 80794 255454 81414 290898
rect 80794 255218 80826 255454
rect 81062 255218 81146 255454
rect 81382 255218 81414 255454
rect 80794 255134 81414 255218
rect 80794 254898 80826 255134
rect 81062 254898 81146 255134
rect 81382 254898 81414 255134
rect 80794 219454 81414 254898
rect 80794 219218 80826 219454
rect 81062 219218 81146 219454
rect 81382 219218 81414 219454
rect 80794 219134 81414 219218
rect 80794 218898 80826 219134
rect 81062 218898 81146 219134
rect 81382 218898 81414 219134
rect 80794 183454 81414 218898
rect 80794 183218 80826 183454
rect 81062 183218 81146 183454
rect 81382 183218 81414 183454
rect 80794 183134 81414 183218
rect 80794 182898 80826 183134
rect 81062 182898 81146 183134
rect 81382 182898 81414 183134
rect 80794 147454 81414 182898
rect 80794 147218 80826 147454
rect 81062 147218 81146 147454
rect 81382 147218 81414 147454
rect 80794 147134 81414 147218
rect 80794 146898 80826 147134
rect 81062 146898 81146 147134
rect 81382 146898 81414 147134
rect 80794 111454 81414 146898
rect 80794 111218 80826 111454
rect 81062 111218 81146 111454
rect 81382 111218 81414 111454
rect 80794 111134 81414 111218
rect 80794 110898 80826 111134
rect 81062 110898 81146 111134
rect 81382 110898 81414 111134
rect 80794 75454 81414 110898
rect 80794 75218 80826 75454
rect 81062 75218 81146 75454
rect 81382 75218 81414 75454
rect 80794 75134 81414 75218
rect 80794 74898 80826 75134
rect 81062 74898 81146 75134
rect 81382 74898 81414 75134
rect 80794 39454 81414 74898
rect 80794 39218 80826 39454
rect 81062 39218 81146 39454
rect 81382 39218 81414 39454
rect 80794 39134 81414 39218
rect 80794 38898 80826 39134
rect 81062 38898 81146 39134
rect 81382 38898 81414 39134
rect 80794 3454 81414 38898
rect 80794 3218 80826 3454
rect 81062 3218 81146 3454
rect 81382 3218 81414 3454
rect 80794 3134 81414 3218
rect 80794 2898 80826 3134
rect 81062 2898 81146 3134
rect 81382 2898 81414 3134
rect 80794 -346 81414 2898
rect 80794 -582 80826 -346
rect 81062 -582 81146 -346
rect 81382 -582 81414 -346
rect 80794 -666 81414 -582
rect 80794 -902 80826 -666
rect 81062 -902 81146 -666
rect 81382 -902 81414 -666
rect 80794 -1894 81414 -902
rect 81954 680614 82574 711002
rect 91954 710598 92574 711590
rect 91954 710362 91986 710598
rect 92222 710362 92306 710598
rect 92542 710362 92574 710598
rect 91954 710278 92574 710362
rect 91954 710042 91986 710278
rect 92222 710042 92306 710278
rect 92542 710042 92574 710278
rect 88234 708678 88854 709670
rect 88234 708442 88266 708678
rect 88502 708442 88586 708678
rect 88822 708442 88854 708678
rect 88234 708358 88854 708442
rect 88234 708122 88266 708358
rect 88502 708122 88586 708358
rect 88822 708122 88854 708358
rect 81954 680378 81986 680614
rect 82222 680378 82306 680614
rect 82542 680378 82574 680614
rect 81954 680294 82574 680378
rect 81954 680058 81986 680294
rect 82222 680058 82306 680294
rect 82542 680058 82574 680294
rect 81954 644614 82574 680058
rect 81954 644378 81986 644614
rect 82222 644378 82306 644614
rect 82542 644378 82574 644614
rect 81954 644294 82574 644378
rect 81954 644058 81986 644294
rect 82222 644058 82306 644294
rect 82542 644058 82574 644294
rect 81954 608614 82574 644058
rect 81954 608378 81986 608614
rect 82222 608378 82306 608614
rect 82542 608378 82574 608614
rect 81954 608294 82574 608378
rect 81954 608058 81986 608294
rect 82222 608058 82306 608294
rect 82542 608058 82574 608294
rect 81954 572614 82574 608058
rect 81954 572378 81986 572614
rect 82222 572378 82306 572614
rect 82542 572378 82574 572614
rect 81954 572294 82574 572378
rect 81954 572058 81986 572294
rect 82222 572058 82306 572294
rect 82542 572058 82574 572294
rect 81954 536614 82574 572058
rect 81954 536378 81986 536614
rect 82222 536378 82306 536614
rect 82542 536378 82574 536614
rect 81954 536294 82574 536378
rect 81954 536058 81986 536294
rect 82222 536058 82306 536294
rect 82542 536058 82574 536294
rect 81954 500614 82574 536058
rect 81954 500378 81986 500614
rect 82222 500378 82306 500614
rect 82542 500378 82574 500614
rect 81954 500294 82574 500378
rect 81954 500058 81986 500294
rect 82222 500058 82306 500294
rect 82542 500058 82574 500294
rect 81954 464614 82574 500058
rect 81954 464378 81986 464614
rect 82222 464378 82306 464614
rect 82542 464378 82574 464614
rect 81954 464294 82574 464378
rect 81954 464058 81986 464294
rect 82222 464058 82306 464294
rect 82542 464058 82574 464294
rect 81954 428614 82574 464058
rect 81954 428378 81986 428614
rect 82222 428378 82306 428614
rect 82542 428378 82574 428614
rect 81954 428294 82574 428378
rect 81954 428058 81986 428294
rect 82222 428058 82306 428294
rect 82542 428058 82574 428294
rect 81954 392614 82574 428058
rect 81954 392378 81986 392614
rect 82222 392378 82306 392614
rect 82542 392378 82574 392614
rect 81954 392294 82574 392378
rect 81954 392058 81986 392294
rect 82222 392058 82306 392294
rect 82542 392058 82574 392294
rect 81954 356614 82574 392058
rect 81954 356378 81986 356614
rect 82222 356378 82306 356614
rect 82542 356378 82574 356614
rect 81954 356294 82574 356378
rect 81954 356058 81986 356294
rect 82222 356058 82306 356294
rect 82542 356058 82574 356294
rect 81954 320614 82574 356058
rect 81954 320378 81986 320614
rect 82222 320378 82306 320614
rect 82542 320378 82574 320614
rect 81954 320294 82574 320378
rect 81954 320058 81986 320294
rect 82222 320058 82306 320294
rect 82542 320058 82574 320294
rect 81954 284614 82574 320058
rect 81954 284378 81986 284614
rect 82222 284378 82306 284614
rect 82542 284378 82574 284614
rect 81954 284294 82574 284378
rect 81954 284058 81986 284294
rect 82222 284058 82306 284294
rect 82542 284058 82574 284294
rect 81954 248614 82574 284058
rect 81954 248378 81986 248614
rect 82222 248378 82306 248614
rect 82542 248378 82574 248614
rect 81954 248294 82574 248378
rect 81954 248058 81986 248294
rect 82222 248058 82306 248294
rect 82542 248058 82574 248294
rect 81954 212614 82574 248058
rect 81954 212378 81986 212614
rect 82222 212378 82306 212614
rect 82542 212378 82574 212614
rect 81954 212294 82574 212378
rect 81954 212058 81986 212294
rect 82222 212058 82306 212294
rect 82542 212058 82574 212294
rect 81954 176614 82574 212058
rect 81954 176378 81986 176614
rect 82222 176378 82306 176614
rect 82542 176378 82574 176614
rect 81954 176294 82574 176378
rect 81954 176058 81986 176294
rect 82222 176058 82306 176294
rect 82542 176058 82574 176294
rect 81954 140614 82574 176058
rect 81954 140378 81986 140614
rect 82222 140378 82306 140614
rect 82542 140378 82574 140614
rect 81954 140294 82574 140378
rect 81954 140058 81986 140294
rect 82222 140058 82306 140294
rect 82542 140058 82574 140294
rect 81954 104614 82574 140058
rect 81954 104378 81986 104614
rect 82222 104378 82306 104614
rect 82542 104378 82574 104614
rect 81954 104294 82574 104378
rect 81954 104058 81986 104294
rect 82222 104058 82306 104294
rect 82542 104058 82574 104294
rect 81954 68614 82574 104058
rect 81954 68378 81986 68614
rect 82222 68378 82306 68614
rect 82542 68378 82574 68614
rect 81954 68294 82574 68378
rect 81954 68058 81986 68294
rect 82222 68058 82306 68294
rect 82542 68058 82574 68294
rect 81954 32614 82574 68058
rect 81954 32378 81986 32614
rect 82222 32378 82306 32614
rect 82542 32378 82574 32614
rect 81954 32294 82574 32378
rect 81954 32058 81986 32294
rect 82222 32058 82306 32294
rect 82542 32058 82574 32294
rect 78234 -5382 78266 -5146
rect 78502 -5382 78586 -5146
rect 78822 -5382 78854 -5146
rect 78234 -5466 78854 -5382
rect 78234 -5702 78266 -5466
rect 78502 -5702 78586 -5466
rect 78822 -5702 78854 -5466
rect 78234 -5734 78854 -5702
rect 71954 -6342 71986 -6106
rect 72222 -6342 72306 -6106
rect 72542 -6342 72574 -6106
rect 71954 -6426 72574 -6342
rect 71954 -6662 71986 -6426
rect 72222 -6662 72306 -6426
rect 72542 -6662 72574 -6426
rect 71954 -7654 72574 -6662
rect 81954 -7066 82574 32058
rect 84514 706758 85134 707750
rect 84514 706522 84546 706758
rect 84782 706522 84866 706758
rect 85102 706522 85134 706758
rect 84514 706438 85134 706522
rect 84514 706202 84546 706438
rect 84782 706202 84866 706438
rect 85102 706202 85134 706438
rect 84514 691174 85134 706202
rect 84514 690938 84546 691174
rect 84782 690938 84866 691174
rect 85102 690938 85134 691174
rect 84514 690854 85134 690938
rect 84514 690618 84546 690854
rect 84782 690618 84866 690854
rect 85102 690618 85134 690854
rect 84514 655174 85134 690618
rect 84514 654938 84546 655174
rect 84782 654938 84866 655174
rect 85102 654938 85134 655174
rect 84514 654854 85134 654938
rect 84514 654618 84546 654854
rect 84782 654618 84866 654854
rect 85102 654618 85134 654854
rect 84514 619174 85134 654618
rect 84514 618938 84546 619174
rect 84782 618938 84866 619174
rect 85102 618938 85134 619174
rect 84514 618854 85134 618938
rect 84514 618618 84546 618854
rect 84782 618618 84866 618854
rect 85102 618618 85134 618854
rect 84514 583174 85134 618618
rect 84514 582938 84546 583174
rect 84782 582938 84866 583174
rect 85102 582938 85134 583174
rect 84514 582854 85134 582938
rect 84514 582618 84546 582854
rect 84782 582618 84866 582854
rect 85102 582618 85134 582854
rect 84514 547174 85134 582618
rect 84514 546938 84546 547174
rect 84782 546938 84866 547174
rect 85102 546938 85134 547174
rect 84514 546854 85134 546938
rect 84514 546618 84546 546854
rect 84782 546618 84866 546854
rect 85102 546618 85134 546854
rect 84514 511174 85134 546618
rect 84514 510938 84546 511174
rect 84782 510938 84866 511174
rect 85102 510938 85134 511174
rect 84514 510854 85134 510938
rect 84514 510618 84546 510854
rect 84782 510618 84866 510854
rect 85102 510618 85134 510854
rect 84514 475174 85134 510618
rect 84514 474938 84546 475174
rect 84782 474938 84866 475174
rect 85102 474938 85134 475174
rect 84514 474854 85134 474938
rect 84514 474618 84546 474854
rect 84782 474618 84866 474854
rect 85102 474618 85134 474854
rect 84514 439174 85134 474618
rect 84514 438938 84546 439174
rect 84782 438938 84866 439174
rect 85102 438938 85134 439174
rect 84514 438854 85134 438938
rect 84514 438618 84546 438854
rect 84782 438618 84866 438854
rect 85102 438618 85134 438854
rect 84514 403174 85134 438618
rect 84514 402938 84546 403174
rect 84782 402938 84866 403174
rect 85102 402938 85134 403174
rect 84514 402854 85134 402938
rect 84514 402618 84546 402854
rect 84782 402618 84866 402854
rect 85102 402618 85134 402854
rect 84514 367174 85134 402618
rect 84514 366938 84546 367174
rect 84782 366938 84866 367174
rect 85102 366938 85134 367174
rect 84514 366854 85134 366938
rect 84514 366618 84546 366854
rect 84782 366618 84866 366854
rect 85102 366618 85134 366854
rect 84514 331174 85134 366618
rect 84514 330938 84546 331174
rect 84782 330938 84866 331174
rect 85102 330938 85134 331174
rect 84514 330854 85134 330938
rect 84514 330618 84546 330854
rect 84782 330618 84866 330854
rect 85102 330618 85134 330854
rect 84514 295174 85134 330618
rect 84514 294938 84546 295174
rect 84782 294938 84866 295174
rect 85102 294938 85134 295174
rect 84514 294854 85134 294938
rect 84514 294618 84546 294854
rect 84782 294618 84866 294854
rect 85102 294618 85134 294854
rect 84514 259174 85134 294618
rect 84514 258938 84546 259174
rect 84782 258938 84866 259174
rect 85102 258938 85134 259174
rect 84514 258854 85134 258938
rect 84514 258618 84546 258854
rect 84782 258618 84866 258854
rect 85102 258618 85134 258854
rect 84514 223174 85134 258618
rect 84514 222938 84546 223174
rect 84782 222938 84866 223174
rect 85102 222938 85134 223174
rect 84514 222854 85134 222938
rect 84514 222618 84546 222854
rect 84782 222618 84866 222854
rect 85102 222618 85134 222854
rect 84514 187174 85134 222618
rect 84514 186938 84546 187174
rect 84782 186938 84866 187174
rect 85102 186938 85134 187174
rect 84514 186854 85134 186938
rect 84514 186618 84546 186854
rect 84782 186618 84866 186854
rect 85102 186618 85134 186854
rect 84514 151174 85134 186618
rect 84514 150938 84546 151174
rect 84782 150938 84866 151174
rect 85102 150938 85134 151174
rect 84514 150854 85134 150938
rect 84514 150618 84546 150854
rect 84782 150618 84866 150854
rect 85102 150618 85134 150854
rect 84514 115174 85134 150618
rect 84514 114938 84546 115174
rect 84782 114938 84866 115174
rect 85102 114938 85134 115174
rect 84514 114854 85134 114938
rect 84514 114618 84546 114854
rect 84782 114618 84866 114854
rect 85102 114618 85134 114854
rect 84514 79174 85134 114618
rect 84514 78938 84546 79174
rect 84782 78938 84866 79174
rect 85102 78938 85134 79174
rect 84514 78854 85134 78938
rect 84514 78618 84546 78854
rect 84782 78618 84866 78854
rect 85102 78618 85134 78854
rect 84514 43174 85134 78618
rect 84514 42938 84546 43174
rect 84782 42938 84866 43174
rect 85102 42938 85134 43174
rect 84514 42854 85134 42938
rect 84514 42618 84546 42854
rect 84782 42618 84866 42854
rect 85102 42618 85134 42854
rect 84514 7174 85134 42618
rect 84514 6938 84546 7174
rect 84782 6938 84866 7174
rect 85102 6938 85134 7174
rect 84514 6854 85134 6938
rect 84514 6618 84546 6854
rect 84782 6618 84866 6854
rect 85102 6618 85134 6854
rect 84514 -2266 85134 6618
rect 84514 -2502 84546 -2266
rect 84782 -2502 84866 -2266
rect 85102 -2502 85134 -2266
rect 84514 -2586 85134 -2502
rect 84514 -2822 84546 -2586
rect 84782 -2822 84866 -2586
rect 85102 -2822 85134 -2586
rect 84514 -3814 85134 -2822
rect 88234 694894 88854 708122
rect 88234 694658 88266 694894
rect 88502 694658 88586 694894
rect 88822 694658 88854 694894
rect 88234 694574 88854 694658
rect 88234 694338 88266 694574
rect 88502 694338 88586 694574
rect 88822 694338 88854 694574
rect 88234 658894 88854 694338
rect 88234 658658 88266 658894
rect 88502 658658 88586 658894
rect 88822 658658 88854 658894
rect 88234 658574 88854 658658
rect 88234 658338 88266 658574
rect 88502 658338 88586 658574
rect 88822 658338 88854 658574
rect 88234 622894 88854 658338
rect 88234 622658 88266 622894
rect 88502 622658 88586 622894
rect 88822 622658 88854 622894
rect 88234 622574 88854 622658
rect 88234 622338 88266 622574
rect 88502 622338 88586 622574
rect 88822 622338 88854 622574
rect 88234 586894 88854 622338
rect 88234 586658 88266 586894
rect 88502 586658 88586 586894
rect 88822 586658 88854 586894
rect 88234 586574 88854 586658
rect 88234 586338 88266 586574
rect 88502 586338 88586 586574
rect 88822 586338 88854 586574
rect 88234 550894 88854 586338
rect 88234 550658 88266 550894
rect 88502 550658 88586 550894
rect 88822 550658 88854 550894
rect 88234 550574 88854 550658
rect 88234 550338 88266 550574
rect 88502 550338 88586 550574
rect 88822 550338 88854 550574
rect 88234 514894 88854 550338
rect 88234 514658 88266 514894
rect 88502 514658 88586 514894
rect 88822 514658 88854 514894
rect 88234 514574 88854 514658
rect 88234 514338 88266 514574
rect 88502 514338 88586 514574
rect 88822 514338 88854 514574
rect 88234 478894 88854 514338
rect 88234 478658 88266 478894
rect 88502 478658 88586 478894
rect 88822 478658 88854 478894
rect 88234 478574 88854 478658
rect 88234 478338 88266 478574
rect 88502 478338 88586 478574
rect 88822 478338 88854 478574
rect 88234 442894 88854 478338
rect 88234 442658 88266 442894
rect 88502 442658 88586 442894
rect 88822 442658 88854 442894
rect 88234 442574 88854 442658
rect 88234 442338 88266 442574
rect 88502 442338 88586 442574
rect 88822 442338 88854 442574
rect 88234 406894 88854 442338
rect 88234 406658 88266 406894
rect 88502 406658 88586 406894
rect 88822 406658 88854 406894
rect 88234 406574 88854 406658
rect 88234 406338 88266 406574
rect 88502 406338 88586 406574
rect 88822 406338 88854 406574
rect 88234 370894 88854 406338
rect 88234 370658 88266 370894
rect 88502 370658 88586 370894
rect 88822 370658 88854 370894
rect 88234 370574 88854 370658
rect 88234 370338 88266 370574
rect 88502 370338 88586 370574
rect 88822 370338 88854 370574
rect 88234 334894 88854 370338
rect 88234 334658 88266 334894
rect 88502 334658 88586 334894
rect 88822 334658 88854 334894
rect 88234 334574 88854 334658
rect 88234 334338 88266 334574
rect 88502 334338 88586 334574
rect 88822 334338 88854 334574
rect 88234 298894 88854 334338
rect 88234 298658 88266 298894
rect 88502 298658 88586 298894
rect 88822 298658 88854 298894
rect 88234 298574 88854 298658
rect 88234 298338 88266 298574
rect 88502 298338 88586 298574
rect 88822 298338 88854 298574
rect 88234 262894 88854 298338
rect 88234 262658 88266 262894
rect 88502 262658 88586 262894
rect 88822 262658 88854 262894
rect 88234 262574 88854 262658
rect 88234 262338 88266 262574
rect 88502 262338 88586 262574
rect 88822 262338 88854 262574
rect 88234 226894 88854 262338
rect 88234 226658 88266 226894
rect 88502 226658 88586 226894
rect 88822 226658 88854 226894
rect 88234 226574 88854 226658
rect 88234 226338 88266 226574
rect 88502 226338 88586 226574
rect 88822 226338 88854 226574
rect 88234 190894 88854 226338
rect 88234 190658 88266 190894
rect 88502 190658 88586 190894
rect 88822 190658 88854 190894
rect 88234 190574 88854 190658
rect 88234 190338 88266 190574
rect 88502 190338 88586 190574
rect 88822 190338 88854 190574
rect 88234 154894 88854 190338
rect 88234 154658 88266 154894
rect 88502 154658 88586 154894
rect 88822 154658 88854 154894
rect 88234 154574 88854 154658
rect 88234 154338 88266 154574
rect 88502 154338 88586 154574
rect 88822 154338 88854 154574
rect 88234 118894 88854 154338
rect 88234 118658 88266 118894
rect 88502 118658 88586 118894
rect 88822 118658 88854 118894
rect 88234 118574 88854 118658
rect 88234 118338 88266 118574
rect 88502 118338 88586 118574
rect 88822 118338 88854 118574
rect 88234 82894 88854 118338
rect 88234 82658 88266 82894
rect 88502 82658 88586 82894
rect 88822 82658 88854 82894
rect 88234 82574 88854 82658
rect 88234 82338 88266 82574
rect 88502 82338 88586 82574
rect 88822 82338 88854 82574
rect 88234 46894 88854 82338
rect 88234 46658 88266 46894
rect 88502 46658 88586 46894
rect 88822 46658 88854 46894
rect 88234 46574 88854 46658
rect 88234 46338 88266 46574
rect 88502 46338 88586 46574
rect 88822 46338 88854 46574
rect 88234 10894 88854 46338
rect 88234 10658 88266 10894
rect 88502 10658 88586 10894
rect 88822 10658 88854 10894
rect 88234 10574 88854 10658
rect 88234 10338 88266 10574
rect 88502 10338 88586 10574
rect 88822 10338 88854 10574
rect 88234 -4186 88854 10338
rect 90794 705798 91414 705830
rect 90794 705562 90826 705798
rect 91062 705562 91146 705798
rect 91382 705562 91414 705798
rect 90794 705478 91414 705562
rect 90794 705242 90826 705478
rect 91062 705242 91146 705478
rect 91382 705242 91414 705478
rect 90794 669454 91414 705242
rect 90794 669218 90826 669454
rect 91062 669218 91146 669454
rect 91382 669218 91414 669454
rect 90794 669134 91414 669218
rect 90794 668898 90826 669134
rect 91062 668898 91146 669134
rect 91382 668898 91414 669134
rect 90794 633454 91414 668898
rect 90794 633218 90826 633454
rect 91062 633218 91146 633454
rect 91382 633218 91414 633454
rect 90794 633134 91414 633218
rect 90794 632898 90826 633134
rect 91062 632898 91146 633134
rect 91382 632898 91414 633134
rect 90794 597454 91414 632898
rect 90794 597218 90826 597454
rect 91062 597218 91146 597454
rect 91382 597218 91414 597454
rect 90794 597134 91414 597218
rect 90794 596898 90826 597134
rect 91062 596898 91146 597134
rect 91382 596898 91414 597134
rect 90794 561454 91414 596898
rect 90794 561218 90826 561454
rect 91062 561218 91146 561454
rect 91382 561218 91414 561454
rect 90794 561134 91414 561218
rect 90794 560898 90826 561134
rect 91062 560898 91146 561134
rect 91382 560898 91414 561134
rect 90794 525454 91414 560898
rect 90794 525218 90826 525454
rect 91062 525218 91146 525454
rect 91382 525218 91414 525454
rect 90794 525134 91414 525218
rect 90794 524898 90826 525134
rect 91062 524898 91146 525134
rect 91382 524898 91414 525134
rect 90794 489454 91414 524898
rect 90794 489218 90826 489454
rect 91062 489218 91146 489454
rect 91382 489218 91414 489454
rect 90794 489134 91414 489218
rect 90794 488898 90826 489134
rect 91062 488898 91146 489134
rect 91382 488898 91414 489134
rect 90794 453454 91414 488898
rect 90794 453218 90826 453454
rect 91062 453218 91146 453454
rect 91382 453218 91414 453454
rect 90794 453134 91414 453218
rect 90794 452898 90826 453134
rect 91062 452898 91146 453134
rect 91382 452898 91414 453134
rect 90794 417454 91414 452898
rect 90794 417218 90826 417454
rect 91062 417218 91146 417454
rect 91382 417218 91414 417454
rect 90794 417134 91414 417218
rect 90794 416898 90826 417134
rect 91062 416898 91146 417134
rect 91382 416898 91414 417134
rect 90794 381454 91414 416898
rect 90794 381218 90826 381454
rect 91062 381218 91146 381454
rect 91382 381218 91414 381454
rect 90794 381134 91414 381218
rect 90794 380898 90826 381134
rect 91062 380898 91146 381134
rect 91382 380898 91414 381134
rect 90794 345454 91414 380898
rect 90794 345218 90826 345454
rect 91062 345218 91146 345454
rect 91382 345218 91414 345454
rect 90794 345134 91414 345218
rect 90794 344898 90826 345134
rect 91062 344898 91146 345134
rect 91382 344898 91414 345134
rect 90794 309454 91414 344898
rect 90794 309218 90826 309454
rect 91062 309218 91146 309454
rect 91382 309218 91414 309454
rect 90794 309134 91414 309218
rect 90794 308898 90826 309134
rect 91062 308898 91146 309134
rect 91382 308898 91414 309134
rect 90794 273454 91414 308898
rect 90794 273218 90826 273454
rect 91062 273218 91146 273454
rect 91382 273218 91414 273454
rect 90794 273134 91414 273218
rect 90794 272898 90826 273134
rect 91062 272898 91146 273134
rect 91382 272898 91414 273134
rect 90794 237454 91414 272898
rect 90794 237218 90826 237454
rect 91062 237218 91146 237454
rect 91382 237218 91414 237454
rect 90794 237134 91414 237218
rect 90794 236898 90826 237134
rect 91062 236898 91146 237134
rect 91382 236898 91414 237134
rect 90794 201454 91414 236898
rect 90794 201218 90826 201454
rect 91062 201218 91146 201454
rect 91382 201218 91414 201454
rect 90794 201134 91414 201218
rect 90794 200898 90826 201134
rect 91062 200898 91146 201134
rect 91382 200898 91414 201134
rect 90794 165454 91414 200898
rect 90794 165218 90826 165454
rect 91062 165218 91146 165454
rect 91382 165218 91414 165454
rect 90794 165134 91414 165218
rect 90794 164898 90826 165134
rect 91062 164898 91146 165134
rect 91382 164898 91414 165134
rect 90794 129454 91414 164898
rect 90794 129218 90826 129454
rect 91062 129218 91146 129454
rect 91382 129218 91414 129454
rect 90794 129134 91414 129218
rect 90794 128898 90826 129134
rect 91062 128898 91146 129134
rect 91382 128898 91414 129134
rect 90794 93454 91414 128898
rect 90794 93218 90826 93454
rect 91062 93218 91146 93454
rect 91382 93218 91414 93454
rect 90794 93134 91414 93218
rect 90794 92898 90826 93134
rect 91062 92898 91146 93134
rect 91382 92898 91414 93134
rect 90794 57454 91414 92898
rect 90794 57218 90826 57454
rect 91062 57218 91146 57454
rect 91382 57218 91414 57454
rect 90794 57134 91414 57218
rect 90794 56898 90826 57134
rect 91062 56898 91146 57134
rect 91382 56898 91414 57134
rect 90794 21454 91414 56898
rect 90794 21218 90826 21454
rect 91062 21218 91146 21454
rect 91382 21218 91414 21454
rect 90794 21134 91414 21218
rect 90794 20898 90826 21134
rect 91062 20898 91146 21134
rect 91382 20898 91414 21134
rect 90794 -1306 91414 20898
rect 90794 -1542 90826 -1306
rect 91062 -1542 91146 -1306
rect 91382 -1542 91414 -1306
rect 90794 -1626 91414 -1542
rect 90794 -1862 90826 -1626
rect 91062 -1862 91146 -1626
rect 91382 -1862 91414 -1626
rect 90794 -1894 91414 -1862
rect 91954 698614 92574 710042
rect 101954 711558 102574 711590
rect 101954 711322 101986 711558
rect 102222 711322 102306 711558
rect 102542 711322 102574 711558
rect 101954 711238 102574 711322
rect 101954 711002 101986 711238
rect 102222 711002 102306 711238
rect 102542 711002 102574 711238
rect 98234 709638 98854 709670
rect 98234 709402 98266 709638
rect 98502 709402 98586 709638
rect 98822 709402 98854 709638
rect 98234 709318 98854 709402
rect 98234 709082 98266 709318
rect 98502 709082 98586 709318
rect 98822 709082 98854 709318
rect 91954 698378 91986 698614
rect 92222 698378 92306 698614
rect 92542 698378 92574 698614
rect 91954 698294 92574 698378
rect 91954 698058 91986 698294
rect 92222 698058 92306 698294
rect 92542 698058 92574 698294
rect 91954 662614 92574 698058
rect 91954 662378 91986 662614
rect 92222 662378 92306 662614
rect 92542 662378 92574 662614
rect 91954 662294 92574 662378
rect 91954 662058 91986 662294
rect 92222 662058 92306 662294
rect 92542 662058 92574 662294
rect 91954 626614 92574 662058
rect 91954 626378 91986 626614
rect 92222 626378 92306 626614
rect 92542 626378 92574 626614
rect 91954 626294 92574 626378
rect 91954 626058 91986 626294
rect 92222 626058 92306 626294
rect 92542 626058 92574 626294
rect 91954 590614 92574 626058
rect 91954 590378 91986 590614
rect 92222 590378 92306 590614
rect 92542 590378 92574 590614
rect 91954 590294 92574 590378
rect 91954 590058 91986 590294
rect 92222 590058 92306 590294
rect 92542 590058 92574 590294
rect 91954 554614 92574 590058
rect 91954 554378 91986 554614
rect 92222 554378 92306 554614
rect 92542 554378 92574 554614
rect 91954 554294 92574 554378
rect 91954 554058 91986 554294
rect 92222 554058 92306 554294
rect 92542 554058 92574 554294
rect 91954 518614 92574 554058
rect 91954 518378 91986 518614
rect 92222 518378 92306 518614
rect 92542 518378 92574 518614
rect 91954 518294 92574 518378
rect 91954 518058 91986 518294
rect 92222 518058 92306 518294
rect 92542 518058 92574 518294
rect 91954 482614 92574 518058
rect 91954 482378 91986 482614
rect 92222 482378 92306 482614
rect 92542 482378 92574 482614
rect 91954 482294 92574 482378
rect 91954 482058 91986 482294
rect 92222 482058 92306 482294
rect 92542 482058 92574 482294
rect 91954 446614 92574 482058
rect 91954 446378 91986 446614
rect 92222 446378 92306 446614
rect 92542 446378 92574 446614
rect 91954 446294 92574 446378
rect 91954 446058 91986 446294
rect 92222 446058 92306 446294
rect 92542 446058 92574 446294
rect 91954 410614 92574 446058
rect 91954 410378 91986 410614
rect 92222 410378 92306 410614
rect 92542 410378 92574 410614
rect 91954 410294 92574 410378
rect 91954 410058 91986 410294
rect 92222 410058 92306 410294
rect 92542 410058 92574 410294
rect 91954 374614 92574 410058
rect 91954 374378 91986 374614
rect 92222 374378 92306 374614
rect 92542 374378 92574 374614
rect 91954 374294 92574 374378
rect 91954 374058 91986 374294
rect 92222 374058 92306 374294
rect 92542 374058 92574 374294
rect 91954 338614 92574 374058
rect 91954 338378 91986 338614
rect 92222 338378 92306 338614
rect 92542 338378 92574 338614
rect 91954 338294 92574 338378
rect 91954 338058 91986 338294
rect 92222 338058 92306 338294
rect 92542 338058 92574 338294
rect 91954 302614 92574 338058
rect 91954 302378 91986 302614
rect 92222 302378 92306 302614
rect 92542 302378 92574 302614
rect 91954 302294 92574 302378
rect 91954 302058 91986 302294
rect 92222 302058 92306 302294
rect 92542 302058 92574 302294
rect 91954 266614 92574 302058
rect 91954 266378 91986 266614
rect 92222 266378 92306 266614
rect 92542 266378 92574 266614
rect 91954 266294 92574 266378
rect 91954 266058 91986 266294
rect 92222 266058 92306 266294
rect 92542 266058 92574 266294
rect 91954 230614 92574 266058
rect 91954 230378 91986 230614
rect 92222 230378 92306 230614
rect 92542 230378 92574 230614
rect 91954 230294 92574 230378
rect 91954 230058 91986 230294
rect 92222 230058 92306 230294
rect 92542 230058 92574 230294
rect 91954 194614 92574 230058
rect 91954 194378 91986 194614
rect 92222 194378 92306 194614
rect 92542 194378 92574 194614
rect 91954 194294 92574 194378
rect 91954 194058 91986 194294
rect 92222 194058 92306 194294
rect 92542 194058 92574 194294
rect 91954 158614 92574 194058
rect 91954 158378 91986 158614
rect 92222 158378 92306 158614
rect 92542 158378 92574 158614
rect 91954 158294 92574 158378
rect 91954 158058 91986 158294
rect 92222 158058 92306 158294
rect 92542 158058 92574 158294
rect 91954 122614 92574 158058
rect 91954 122378 91986 122614
rect 92222 122378 92306 122614
rect 92542 122378 92574 122614
rect 91954 122294 92574 122378
rect 91954 122058 91986 122294
rect 92222 122058 92306 122294
rect 92542 122058 92574 122294
rect 91954 86614 92574 122058
rect 91954 86378 91986 86614
rect 92222 86378 92306 86614
rect 92542 86378 92574 86614
rect 91954 86294 92574 86378
rect 91954 86058 91986 86294
rect 92222 86058 92306 86294
rect 92542 86058 92574 86294
rect 91954 50614 92574 86058
rect 91954 50378 91986 50614
rect 92222 50378 92306 50614
rect 92542 50378 92574 50614
rect 91954 50294 92574 50378
rect 91954 50058 91986 50294
rect 92222 50058 92306 50294
rect 92542 50058 92574 50294
rect 91954 14614 92574 50058
rect 91954 14378 91986 14614
rect 92222 14378 92306 14614
rect 92542 14378 92574 14614
rect 91954 14294 92574 14378
rect 91954 14058 91986 14294
rect 92222 14058 92306 14294
rect 92542 14058 92574 14294
rect 88234 -4422 88266 -4186
rect 88502 -4422 88586 -4186
rect 88822 -4422 88854 -4186
rect 88234 -4506 88854 -4422
rect 88234 -4742 88266 -4506
rect 88502 -4742 88586 -4506
rect 88822 -4742 88854 -4506
rect 88234 -5734 88854 -4742
rect 81954 -7302 81986 -7066
rect 82222 -7302 82306 -7066
rect 82542 -7302 82574 -7066
rect 81954 -7386 82574 -7302
rect 81954 -7622 81986 -7386
rect 82222 -7622 82306 -7386
rect 82542 -7622 82574 -7386
rect 81954 -7654 82574 -7622
rect 91954 -6106 92574 14058
rect 94514 707718 95134 707750
rect 94514 707482 94546 707718
rect 94782 707482 94866 707718
rect 95102 707482 95134 707718
rect 94514 707398 95134 707482
rect 94514 707162 94546 707398
rect 94782 707162 94866 707398
rect 95102 707162 95134 707398
rect 94514 673174 95134 707162
rect 94514 672938 94546 673174
rect 94782 672938 94866 673174
rect 95102 672938 95134 673174
rect 94514 672854 95134 672938
rect 94514 672618 94546 672854
rect 94782 672618 94866 672854
rect 95102 672618 95134 672854
rect 94514 637174 95134 672618
rect 94514 636938 94546 637174
rect 94782 636938 94866 637174
rect 95102 636938 95134 637174
rect 94514 636854 95134 636938
rect 94514 636618 94546 636854
rect 94782 636618 94866 636854
rect 95102 636618 95134 636854
rect 94514 601174 95134 636618
rect 94514 600938 94546 601174
rect 94782 600938 94866 601174
rect 95102 600938 95134 601174
rect 94514 600854 95134 600938
rect 94514 600618 94546 600854
rect 94782 600618 94866 600854
rect 95102 600618 95134 600854
rect 94514 565174 95134 600618
rect 94514 564938 94546 565174
rect 94782 564938 94866 565174
rect 95102 564938 95134 565174
rect 94514 564854 95134 564938
rect 94514 564618 94546 564854
rect 94782 564618 94866 564854
rect 95102 564618 95134 564854
rect 94514 529174 95134 564618
rect 94514 528938 94546 529174
rect 94782 528938 94866 529174
rect 95102 528938 95134 529174
rect 94514 528854 95134 528938
rect 94514 528618 94546 528854
rect 94782 528618 94866 528854
rect 95102 528618 95134 528854
rect 94514 493174 95134 528618
rect 94514 492938 94546 493174
rect 94782 492938 94866 493174
rect 95102 492938 95134 493174
rect 94514 492854 95134 492938
rect 94514 492618 94546 492854
rect 94782 492618 94866 492854
rect 95102 492618 95134 492854
rect 94514 457174 95134 492618
rect 94514 456938 94546 457174
rect 94782 456938 94866 457174
rect 95102 456938 95134 457174
rect 94514 456854 95134 456938
rect 94514 456618 94546 456854
rect 94782 456618 94866 456854
rect 95102 456618 95134 456854
rect 94514 421174 95134 456618
rect 94514 420938 94546 421174
rect 94782 420938 94866 421174
rect 95102 420938 95134 421174
rect 94514 420854 95134 420938
rect 94514 420618 94546 420854
rect 94782 420618 94866 420854
rect 95102 420618 95134 420854
rect 94514 385174 95134 420618
rect 94514 384938 94546 385174
rect 94782 384938 94866 385174
rect 95102 384938 95134 385174
rect 94514 384854 95134 384938
rect 94514 384618 94546 384854
rect 94782 384618 94866 384854
rect 95102 384618 95134 384854
rect 94514 349174 95134 384618
rect 94514 348938 94546 349174
rect 94782 348938 94866 349174
rect 95102 348938 95134 349174
rect 94514 348854 95134 348938
rect 94514 348618 94546 348854
rect 94782 348618 94866 348854
rect 95102 348618 95134 348854
rect 94514 313174 95134 348618
rect 94514 312938 94546 313174
rect 94782 312938 94866 313174
rect 95102 312938 95134 313174
rect 94514 312854 95134 312938
rect 94514 312618 94546 312854
rect 94782 312618 94866 312854
rect 95102 312618 95134 312854
rect 94514 277174 95134 312618
rect 94514 276938 94546 277174
rect 94782 276938 94866 277174
rect 95102 276938 95134 277174
rect 94514 276854 95134 276938
rect 94514 276618 94546 276854
rect 94782 276618 94866 276854
rect 95102 276618 95134 276854
rect 94514 241174 95134 276618
rect 94514 240938 94546 241174
rect 94782 240938 94866 241174
rect 95102 240938 95134 241174
rect 94514 240854 95134 240938
rect 94514 240618 94546 240854
rect 94782 240618 94866 240854
rect 95102 240618 95134 240854
rect 94514 205174 95134 240618
rect 94514 204938 94546 205174
rect 94782 204938 94866 205174
rect 95102 204938 95134 205174
rect 94514 204854 95134 204938
rect 94514 204618 94546 204854
rect 94782 204618 94866 204854
rect 95102 204618 95134 204854
rect 94514 169174 95134 204618
rect 94514 168938 94546 169174
rect 94782 168938 94866 169174
rect 95102 168938 95134 169174
rect 94514 168854 95134 168938
rect 94514 168618 94546 168854
rect 94782 168618 94866 168854
rect 95102 168618 95134 168854
rect 94514 133174 95134 168618
rect 94514 132938 94546 133174
rect 94782 132938 94866 133174
rect 95102 132938 95134 133174
rect 94514 132854 95134 132938
rect 94514 132618 94546 132854
rect 94782 132618 94866 132854
rect 95102 132618 95134 132854
rect 94514 97174 95134 132618
rect 94514 96938 94546 97174
rect 94782 96938 94866 97174
rect 95102 96938 95134 97174
rect 94514 96854 95134 96938
rect 94514 96618 94546 96854
rect 94782 96618 94866 96854
rect 95102 96618 95134 96854
rect 94514 61174 95134 96618
rect 94514 60938 94546 61174
rect 94782 60938 94866 61174
rect 95102 60938 95134 61174
rect 94514 60854 95134 60938
rect 94514 60618 94546 60854
rect 94782 60618 94866 60854
rect 95102 60618 95134 60854
rect 94514 25174 95134 60618
rect 94514 24938 94546 25174
rect 94782 24938 94866 25174
rect 95102 24938 95134 25174
rect 94514 24854 95134 24938
rect 94514 24618 94546 24854
rect 94782 24618 94866 24854
rect 95102 24618 95134 24854
rect 94514 -3226 95134 24618
rect 94514 -3462 94546 -3226
rect 94782 -3462 94866 -3226
rect 95102 -3462 95134 -3226
rect 94514 -3546 95134 -3462
rect 94514 -3782 94546 -3546
rect 94782 -3782 94866 -3546
rect 95102 -3782 95134 -3546
rect 94514 -3814 95134 -3782
rect 98234 676894 98854 709082
rect 98234 676658 98266 676894
rect 98502 676658 98586 676894
rect 98822 676658 98854 676894
rect 98234 676574 98854 676658
rect 98234 676338 98266 676574
rect 98502 676338 98586 676574
rect 98822 676338 98854 676574
rect 98234 640894 98854 676338
rect 98234 640658 98266 640894
rect 98502 640658 98586 640894
rect 98822 640658 98854 640894
rect 98234 640574 98854 640658
rect 98234 640338 98266 640574
rect 98502 640338 98586 640574
rect 98822 640338 98854 640574
rect 98234 604894 98854 640338
rect 98234 604658 98266 604894
rect 98502 604658 98586 604894
rect 98822 604658 98854 604894
rect 98234 604574 98854 604658
rect 98234 604338 98266 604574
rect 98502 604338 98586 604574
rect 98822 604338 98854 604574
rect 98234 568894 98854 604338
rect 98234 568658 98266 568894
rect 98502 568658 98586 568894
rect 98822 568658 98854 568894
rect 98234 568574 98854 568658
rect 98234 568338 98266 568574
rect 98502 568338 98586 568574
rect 98822 568338 98854 568574
rect 98234 532894 98854 568338
rect 98234 532658 98266 532894
rect 98502 532658 98586 532894
rect 98822 532658 98854 532894
rect 98234 532574 98854 532658
rect 98234 532338 98266 532574
rect 98502 532338 98586 532574
rect 98822 532338 98854 532574
rect 98234 496894 98854 532338
rect 98234 496658 98266 496894
rect 98502 496658 98586 496894
rect 98822 496658 98854 496894
rect 98234 496574 98854 496658
rect 98234 496338 98266 496574
rect 98502 496338 98586 496574
rect 98822 496338 98854 496574
rect 98234 460894 98854 496338
rect 98234 460658 98266 460894
rect 98502 460658 98586 460894
rect 98822 460658 98854 460894
rect 98234 460574 98854 460658
rect 98234 460338 98266 460574
rect 98502 460338 98586 460574
rect 98822 460338 98854 460574
rect 98234 424894 98854 460338
rect 98234 424658 98266 424894
rect 98502 424658 98586 424894
rect 98822 424658 98854 424894
rect 98234 424574 98854 424658
rect 98234 424338 98266 424574
rect 98502 424338 98586 424574
rect 98822 424338 98854 424574
rect 98234 388894 98854 424338
rect 98234 388658 98266 388894
rect 98502 388658 98586 388894
rect 98822 388658 98854 388894
rect 98234 388574 98854 388658
rect 98234 388338 98266 388574
rect 98502 388338 98586 388574
rect 98822 388338 98854 388574
rect 98234 352894 98854 388338
rect 98234 352658 98266 352894
rect 98502 352658 98586 352894
rect 98822 352658 98854 352894
rect 98234 352574 98854 352658
rect 98234 352338 98266 352574
rect 98502 352338 98586 352574
rect 98822 352338 98854 352574
rect 98234 316894 98854 352338
rect 98234 316658 98266 316894
rect 98502 316658 98586 316894
rect 98822 316658 98854 316894
rect 98234 316574 98854 316658
rect 98234 316338 98266 316574
rect 98502 316338 98586 316574
rect 98822 316338 98854 316574
rect 98234 280894 98854 316338
rect 98234 280658 98266 280894
rect 98502 280658 98586 280894
rect 98822 280658 98854 280894
rect 98234 280574 98854 280658
rect 98234 280338 98266 280574
rect 98502 280338 98586 280574
rect 98822 280338 98854 280574
rect 98234 244894 98854 280338
rect 98234 244658 98266 244894
rect 98502 244658 98586 244894
rect 98822 244658 98854 244894
rect 98234 244574 98854 244658
rect 98234 244338 98266 244574
rect 98502 244338 98586 244574
rect 98822 244338 98854 244574
rect 98234 208894 98854 244338
rect 98234 208658 98266 208894
rect 98502 208658 98586 208894
rect 98822 208658 98854 208894
rect 98234 208574 98854 208658
rect 98234 208338 98266 208574
rect 98502 208338 98586 208574
rect 98822 208338 98854 208574
rect 98234 172894 98854 208338
rect 98234 172658 98266 172894
rect 98502 172658 98586 172894
rect 98822 172658 98854 172894
rect 98234 172574 98854 172658
rect 98234 172338 98266 172574
rect 98502 172338 98586 172574
rect 98822 172338 98854 172574
rect 98234 136894 98854 172338
rect 98234 136658 98266 136894
rect 98502 136658 98586 136894
rect 98822 136658 98854 136894
rect 98234 136574 98854 136658
rect 98234 136338 98266 136574
rect 98502 136338 98586 136574
rect 98822 136338 98854 136574
rect 98234 100894 98854 136338
rect 98234 100658 98266 100894
rect 98502 100658 98586 100894
rect 98822 100658 98854 100894
rect 98234 100574 98854 100658
rect 98234 100338 98266 100574
rect 98502 100338 98586 100574
rect 98822 100338 98854 100574
rect 98234 64894 98854 100338
rect 98234 64658 98266 64894
rect 98502 64658 98586 64894
rect 98822 64658 98854 64894
rect 98234 64574 98854 64658
rect 98234 64338 98266 64574
rect 98502 64338 98586 64574
rect 98822 64338 98854 64574
rect 98234 28894 98854 64338
rect 98234 28658 98266 28894
rect 98502 28658 98586 28894
rect 98822 28658 98854 28894
rect 98234 28574 98854 28658
rect 98234 28338 98266 28574
rect 98502 28338 98586 28574
rect 98822 28338 98854 28574
rect 98234 -5146 98854 28338
rect 100794 704838 101414 705830
rect 100794 704602 100826 704838
rect 101062 704602 101146 704838
rect 101382 704602 101414 704838
rect 100794 704518 101414 704602
rect 100794 704282 100826 704518
rect 101062 704282 101146 704518
rect 101382 704282 101414 704518
rect 100794 687454 101414 704282
rect 100794 687218 100826 687454
rect 101062 687218 101146 687454
rect 101382 687218 101414 687454
rect 100794 687134 101414 687218
rect 100794 686898 100826 687134
rect 101062 686898 101146 687134
rect 101382 686898 101414 687134
rect 100794 651454 101414 686898
rect 100794 651218 100826 651454
rect 101062 651218 101146 651454
rect 101382 651218 101414 651454
rect 100794 651134 101414 651218
rect 100794 650898 100826 651134
rect 101062 650898 101146 651134
rect 101382 650898 101414 651134
rect 100794 615454 101414 650898
rect 100794 615218 100826 615454
rect 101062 615218 101146 615454
rect 101382 615218 101414 615454
rect 100794 615134 101414 615218
rect 100794 614898 100826 615134
rect 101062 614898 101146 615134
rect 101382 614898 101414 615134
rect 100794 579454 101414 614898
rect 100794 579218 100826 579454
rect 101062 579218 101146 579454
rect 101382 579218 101414 579454
rect 100794 579134 101414 579218
rect 100794 578898 100826 579134
rect 101062 578898 101146 579134
rect 101382 578898 101414 579134
rect 100794 543454 101414 578898
rect 100794 543218 100826 543454
rect 101062 543218 101146 543454
rect 101382 543218 101414 543454
rect 100794 543134 101414 543218
rect 100794 542898 100826 543134
rect 101062 542898 101146 543134
rect 101382 542898 101414 543134
rect 100794 507454 101414 542898
rect 100794 507218 100826 507454
rect 101062 507218 101146 507454
rect 101382 507218 101414 507454
rect 100794 507134 101414 507218
rect 100794 506898 100826 507134
rect 101062 506898 101146 507134
rect 101382 506898 101414 507134
rect 100794 471454 101414 506898
rect 100794 471218 100826 471454
rect 101062 471218 101146 471454
rect 101382 471218 101414 471454
rect 100794 471134 101414 471218
rect 100794 470898 100826 471134
rect 101062 470898 101146 471134
rect 101382 470898 101414 471134
rect 100794 435454 101414 470898
rect 100794 435218 100826 435454
rect 101062 435218 101146 435454
rect 101382 435218 101414 435454
rect 100794 435134 101414 435218
rect 100794 434898 100826 435134
rect 101062 434898 101146 435134
rect 101382 434898 101414 435134
rect 100794 399454 101414 434898
rect 100794 399218 100826 399454
rect 101062 399218 101146 399454
rect 101382 399218 101414 399454
rect 100794 399134 101414 399218
rect 100794 398898 100826 399134
rect 101062 398898 101146 399134
rect 101382 398898 101414 399134
rect 100794 363454 101414 398898
rect 100794 363218 100826 363454
rect 101062 363218 101146 363454
rect 101382 363218 101414 363454
rect 100794 363134 101414 363218
rect 100794 362898 100826 363134
rect 101062 362898 101146 363134
rect 101382 362898 101414 363134
rect 100794 327454 101414 362898
rect 100794 327218 100826 327454
rect 101062 327218 101146 327454
rect 101382 327218 101414 327454
rect 100794 327134 101414 327218
rect 100794 326898 100826 327134
rect 101062 326898 101146 327134
rect 101382 326898 101414 327134
rect 100794 291454 101414 326898
rect 100794 291218 100826 291454
rect 101062 291218 101146 291454
rect 101382 291218 101414 291454
rect 100794 291134 101414 291218
rect 100794 290898 100826 291134
rect 101062 290898 101146 291134
rect 101382 290898 101414 291134
rect 100794 255454 101414 290898
rect 100794 255218 100826 255454
rect 101062 255218 101146 255454
rect 101382 255218 101414 255454
rect 100794 255134 101414 255218
rect 100794 254898 100826 255134
rect 101062 254898 101146 255134
rect 101382 254898 101414 255134
rect 100794 219454 101414 254898
rect 100794 219218 100826 219454
rect 101062 219218 101146 219454
rect 101382 219218 101414 219454
rect 100794 219134 101414 219218
rect 100794 218898 100826 219134
rect 101062 218898 101146 219134
rect 101382 218898 101414 219134
rect 100794 183454 101414 218898
rect 100794 183218 100826 183454
rect 101062 183218 101146 183454
rect 101382 183218 101414 183454
rect 100794 183134 101414 183218
rect 100794 182898 100826 183134
rect 101062 182898 101146 183134
rect 101382 182898 101414 183134
rect 100794 147454 101414 182898
rect 100794 147218 100826 147454
rect 101062 147218 101146 147454
rect 101382 147218 101414 147454
rect 100794 147134 101414 147218
rect 100794 146898 100826 147134
rect 101062 146898 101146 147134
rect 101382 146898 101414 147134
rect 100794 111454 101414 146898
rect 100794 111218 100826 111454
rect 101062 111218 101146 111454
rect 101382 111218 101414 111454
rect 100794 111134 101414 111218
rect 100794 110898 100826 111134
rect 101062 110898 101146 111134
rect 101382 110898 101414 111134
rect 100794 75454 101414 110898
rect 100794 75218 100826 75454
rect 101062 75218 101146 75454
rect 101382 75218 101414 75454
rect 100794 75134 101414 75218
rect 100794 74898 100826 75134
rect 101062 74898 101146 75134
rect 101382 74898 101414 75134
rect 100794 39454 101414 74898
rect 100794 39218 100826 39454
rect 101062 39218 101146 39454
rect 101382 39218 101414 39454
rect 100794 39134 101414 39218
rect 100794 38898 100826 39134
rect 101062 38898 101146 39134
rect 101382 38898 101414 39134
rect 100794 3454 101414 38898
rect 100794 3218 100826 3454
rect 101062 3218 101146 3454
rect 101382 3218 101414 3454
rect 100794 3134 101414 3218
rect 100794 2898 100826 3134
rect 101062 2898 101146 3134
rect 101382 2898 101414 3134
rect 100794 -346 101414 2898
rect 100794 -582 100826 -346
rect 101062 -582 101146 -346
rect 101382 -582 101414 -346
rect 100794 -666 101414 -582
rect 100794 -902 100826 -666
rect 101062 -902 101146 -666
rect 101382 -902 101414 -666
rect 100794 -1894 101414 -902
rect 101954 680614 102574 711002
rect 111954 710598 112574 711590
rect 111954 710362 111986 710598
rect 112222 710362 112306 710598
rect 112542 710362 112574 710598
rect 111954 710278 112574 710362
rect 111954 710042 111986 710278
rect 112222 710042 112306 710278
rect 112542 710042 112574 710278
rect 108234 708678 108854 709670
rect 108234 708442 108266 708678
rect 108502 708442 108586 708678
rect 108822 708442 108854 708678
rect 108234 708358 108854 708442
rect 108234 708122 108266 708358
rect 108502 708122 108586 708358
rect 108822 708122 108854 708358
rect 101954 680378 101986 680614
rect 102222 680378 102306 680614
rect 102542 680378 102574 680614
rect 101954 680294 102574 680378
rect 101954 680058 101986 680294
rect 102222 680058 102306 680294
rect 102542 680058 102574 680294
rect 101954 644614 102574 680058
rect 101954 644378 101986 644614
rect 102222 644378 102306 644614
rect 102542 644378 102574 644614
rect 101954 644294 102574 644378
rect 101954 644058 101986 644294
rect 102222 644058 102306 644294
rect 102542 644058 102574 644294
rect 101954 608614 102574 644058
rect 101954 608378 101986 608614
rect 102222 608378 102306 608614
rect 102542 608378 102574 608614
rect 101954 608294 102574 608378
rect 101954 608058 101986 608294
rect 102222 608058 102306 608294
rect 102542 608058 102574 608294
rect 101954 572614 102574 608058
rect 101954 572378 101986 572614
rect 102222 572378 102306 572614
rect 102542 572378 102574 572614
rect 101954 572294 102574 572378
rect 101954 572058 101986 572294
rect 102222 572058 102306 572294
rect 102542 572058 102574 572294
rect 101954 536614 102574 572058
rect 101954 536378 101986 536614
rect 102222 536378 102306 536614
rect 102542 536378 102574 536614
rect 101954 536294 102574 536378
rect 101954 536058 101986 536294
rect 102222 536058 102306 536294
rect 102542 536058 102574 536294
rect 101954 500614 102574 536058
rect 101954 500378 101986 500614
rect 102222 500378 102306 500614
rect 102542 500378 102574 500614
rect 101954 500294 102574 500378
rect 101954 500058 101986 500294
rect 102222 500058 102306 500294
rect 102542 500058 102574 500294
rect 101954 464614 102574 500058
rect 101954 464378 101986 464614
rect 102222 464378 102306 464614
rect 102542 464378 102574 464614
rect 101954 464294 102574 464378
rect 101954 464058 101986 464294
rect 102222 464058 102306 464294
rect 102542 464058 102574 464294
rect 101954 428614 102574 464058
rect 101954 428378 101986 428614
rect 102222 428378 102306 428614
rect 102542 428378 102574 428614
rect 101954 428294 102574 428378
rect 101954 428058 101986 428294
rect 102222 428058 102306 428294
rect 102542 428058 102574 428294
rect 101954 392614 102574 428058
rect 101954 392378 101986 392614
rect 102222 392378 102306 392614
rect 102542 392378 102574 392614
rect 101954 392294 102574 392378
rect 101954 392058 101986 392294
rect 102222 392058 102306 392294
rect 102542 392058 102574 392294
rect 101954 356614 102574 392058
rect 101954 356378 101986 356614
rect 102222 356378 102306 356614
rect 102542 356378 102574 356614
rect 101954 356294 102574 356378
rect 101954 356058 101986 356294
rect 102222 356058 102306 356294
rect 102542 356058 102574 356294
rect 101954 320614 102574 356058
rect 101954 320378 101986 320614
rect 102222 320378 102306 320614
rect 102542 320378 102574 320614
rect 101954 320294 102574 320378
rect 101954 320058 101986 320294
rect 102222 320058 102306 320294
rect 102542 320058 102574 320294
rect 101954 284614 102574 320058
rect 101954 284378 101986 284614
rect 102222 284378 102306 284614
rect 102542 284378 102574 284614
rect 101954 284294 102574 284378
rect 101954 284058 101986 284294
rect 102222 284058 102306 284294
rect 102542 284058 102574 284294
rect 101954 248614 102574 284058
rect 101954 248378 101986 248614
rect 102222 248378 102306 248614
rect 102542 248378 102574 248614
rect 101954 248294 102574 248378
rect 101954 248058 101986 248294
rect 102222 248058 102306 248294
rect 102542 248058 102574 248294
rect 101954 212614 102574 248058
rect 101954 212378 101986 212614
rect 102222 212378 102306 212614
rect 102542 212378 102574 212614
rect 101954 212294 102574 212378
rect 101954 212058 101986 212294
rect 102222 212058 102306 212294
rect 102542 212058 102574 212294
rect 101954 176614 102574 212058
rect 101954 176378 101986 176614
rect 102222 176378 102306 176614
rect 102542 176378 102574 176614
rect 101954 176294 102574 176378
rect 101954 176058 101986 176294
rect 102222 176058 102306 176294
rect 102542 176058 102574 176294
rect 101954 140614 102574 176058
rect 101954 140378 101986 140614
rect 102222 140378 102306 140614
rect 102542 140378 102574 140614
rect 101954 140294 102574 140378
rect 101954 140058 101986 140294
rect 102222 140058 102306 140294
rect 102542 140058 102574 140294
rect 101954 104614 102574 140058
rect 101954 104378 101986 104614
rect 102222 104378 102306 104614
rect 102542 104378 102574 104614
rect 101954 104294 102574 104378
rect 101954 104058 101986 104294
rect 102222 104058 102306 104294
rect 102542 104058 102574 104294
rect 101954 68614 102574 104058
rect 101954 68378 101986 68614
rect 102222 68378 102306 68614
rect 102542 68378 102574 68614
rect 101954 68294 102574 68378
rect 101954 68058 101986 68294
rect 102222 68058 102306 68294
rect 102542 68058 102574 68294
rect 101954 32614 102574 68058
rect 101954 32378 101986 32614
rect 102222 32378 102306 32614
rect 102542 32378 102574 32614
rect 101954 32294 102574 32378
rect 101954 32058 101986 32294
rect 102222 32058 102306 32294
rect 102542 32058 102574 32294
rect 98234 -5382 98266 -5146
rect 98502 -5382 98586 -5146
rect 98822 -5382 98854 -5146
rect 98234 -5466 98854 -5382
rect 98234 -5702 98266 -5466
rect 98502 -5702 98586 -5466
rect 98822 -5702 98854 -5466
rect 98234 -5734 98854 -5702
rect 91954 -6342 91986 -6106
rect 92222 -6342 92306 -6106
rect 92542 -6342 92574 -6106
rect 91954 -6426 92574 -6342
rect 91954 -6662 91986 -6426
rect 92222 -6662 92306 -6426
rect 92542 -6662 92574 -6426
rect 91954 -7654 92574 -6662
rect 101954 -7066 102574 32058
rect 104514 706758 105134 707750
rect 104514 706522 104546 706758
rect 104782 706522 104866 706758
rect 105102 706522 105134 706758
rect 104514 706438 105134 706522
rect 104514 706202 104546 706438
rect 104782 706202 104866 706438
rect 105102 706202 105134 706438
rect 104514 691174 105134 706202
rect 104514 690938 104546 691174
rect 104782 690938 104866 691174
rect 105102 690938 105134 691174
rect 104514 690854 105134 690938
rect 104514 690618 104546 690854
rect 104782 690618 104866 690854
rect 105102 690618 105134 690854
rect 104514 655174 105134 690618
rect 104514 654938 104546 655174
rect 104782 654938 104866 655174
rect 105102 654938 105134 655174
rect 104514 654854 105134 654938
rect 104514 654618 104546 654854
rect 104782 654618 104866 654854
rect 105102 654618 105134 654854
rect 104514 619174 105134 654618
rect 104514 618938 104546 619174
rect 104782 618938 104866 619174
rect 105102 618938 105134 619174
rect 104514 618854 105134 618938
rect 104514 618618 104546 618854
rect 104782 618618 104866 618854
rect 105102 618618 105134 618854
rect 104514 583174 105134 618618
rect 104514 582938 104546 583174
rect 104782 582938 104866 583174
rect 105102 582938 105134 583174
rect 104514 582854 105134 582938
rect 104514 582618 104546 582854
rect 104782 582618 104866 582854
rect 105102 582618 105134 582854
rect 104514 547174 105134 582618
rect 104514 546938 104546 547174
rect 104782 546938 104866 547174
rect 105102 546938 105134 547174
rect 104514 546854 105134 546938
rect 104514 546618 104546 546854
rect 104782 546618 104866 546854
rect 105102 546618 105134 546854
rect 104514 511174 105134 546618
rect 104514 510938 104546 511174
rect 104782 510938 104866 511174
rect 105102 510938 105134 511174
rect 104514 510854 105134 510938
rect 104514 510618 104546 510854
rect 104782 510618 104866 510854
rect 105102 510618 105134 510854
rect 104514 475174 105134 510618
rect 104514 474938 104546 475174
rect 104782 474938 104866 475174
rect 105102 474938 105134 475174
rect 104514 474854 105134 474938
rect 104514 474618 104546 474854
rect 104782 474618 104866 474854
rect 105102 474618 105134 474854
rect 104514 439174 105134 474618
rect 104514 438938 104546 439174
rect 104782 438938 104866 439174
rect 105102 438938 105134 439174
rect 104514 438854 105134 438938
rect 104514 438618 104546 438854
rect 104782 438618 104866 438854
rect 105102 438618 105134 438854
rect 104514 403174 105134 438618
rect 104514 402938 104546 403174
rect 104782 402938 104866 403174
rect 105102 402938 105134 403174
rect 104514 402854 105134 402938
rect 104514 402618 104546 402854
rect 104782 402618 104866 402854
rect 105102 402618 105134 402854
rect 104514 367174 105134 402618
rect 104514 366938 104546 367174
rect 104782 366938 104866 367174
rect 105102 366938 105134 367174
rect 104514 366854 105134 366938
rect 104514 366618 104546 366854
rect 104782 366618 104866 366854
rect 105102 366618 105134 366854
rect 104514 331174 105134 366618
rect 104514 330938 104546 331174
rect 104782 330938 104866 331174
rect 105102 330938 105134 331174
rect 104514 330854 105134 330938
rect 104514 330618 104546 330854
rect 104782 330618 104866 330854
rect 105102 330618 105134 330854
rect 104514 295174 105134 330618
rect 104514 294938 104546 295174
rect 104782 294938 104866 295174
rect 105102 294938 105134 295174
rect 104514 294854 105134 294938
rect 104514 294618 104546 294854
rect 104782 294618 104866 294854
rect 105102 294618 105134 294854
rect 104514 259174 105134 294618
rect 104514 258938 104546 259174
rect 104782 258938 104866 259174
rect 105102 258938 105134 259174
rect 104514 258854 105134 258938
rect 104514 258618 104546 258854
rect 104782 258618 104866 258854
rect 105102 258618 105134 258854
rect 104514 223174 105134 258618
rect 104514 222938 104546 223174
rect 104782 222938 104866 223174
rect 105102 222938 105134 223174
rect 104514 222854 105134 222938
rect 104514 222618 104546 222854
rect 104782 222618 104866 222854
rect 105102 222618 105134 222854
rect 104514 187174 105134 222618
rect 104514 186938 104546 187174
rect 104782 186938 104866 187174
rect 105102 186938 105134 187174
rect 104514 186854 105134 186938
rect 104514 186618 104546 186854
rect 104782 186618 104866 186854
rect 105102 186618 105134 186854
rect 104514 151174 105134 186618
rect 104514 150938 104546 151174
rect 104782 150938 104866 151174
rect 105102 150938 105134 151174
rect 104514 150854 105134 150938
rect 104514 150618 104546 150854
rect 104782 150618 104866 150854
rect 105102 150618 105134 150854
rect 104514 115174 105134 150618
rect 104514 114938 104546 115174
rect 104782 114938 104866 115174
rect 105102 114938 105134 115174
rect 104514 114854 105134 114938
rect 104514 114618 104546 114854
rect 104782 114618 104866 114854
rect 105102 114618 105134 114854
rect 104514 79174 105134 114618
rect 104514 78938 104546 79174
rect 104782 78938 104866 79174
rect 105102 78938 105134 79174
rect 104514 78854 105134 78938
rect 104514 78618 104546 78854
rect 104782 78618 104866 78854
rect 105102 78618 105134 78854
rect 104514 43174 105134 78618
rect 104514 42938 104546 43174
rect 104782 42938 104866 43174
rect 105102 42938 105134 43174
rect 104514 42854 105134 42938
rect 104514 42618 104546 42854
rect 104782 42618 104866 42854
rect 105102 42618 105134 42854
rect 104514 7174 105134 42618
rect 104514 6938 104546 7174
rect 104782 6938 104866 7174
rect 105102 6938 105134 7174
rect 104514 6854 105134 6938
rect 104514 6618 104546 6854
rect 104782 6618 104866 6854
rect 105102 6618 105134 6854
rect 104514 -2266 105134 6618
rect 104514 -2502 104546 -2266
rect 104782 -2502 104866 -2266
rect 105102 -2502 105134 -2266
rect 104514 -2586 105134 -2502
rect 104514 -2822 104546 -2586
rect 104782 -2822 104866 -2586
rect 105102 -2822 105134 -2586
rect 104514 -3814 105134 -2822
rect 108234 694894 108854 708122
rect 108234 694658 108266 694894
rect 108502 694658 108586 694894
rect 108822 694658 108854 694894
rect 108234 694574 108854 694658
rect 108234 694338 108266 694574
rect 108502 694338 108586 694574
rect 108822 694338 108854 694574
rect 108234 658894 108854 694338
rect 108234 658658 108266 658894
rect 108502 658658 108586 658894
rect 108822 658658 108854 658894
rect 108234 658574 108854 658658
rect 108234 658338 108266 658574
rect 108502 658338 108586 658574
rect 108822 658338 108854 658574
rect 108234 622894 108854 658338
rect 108234 622658 108266 622894
rect 108502 622658 108586 622894
rect 108822 622658 108854 622894
rect 108234 622574 108854 622658
rect 108234 622338 108266 622574
rect 108502 622338 108586 622574
rect 108822 622338 108854 622574
rect 108234 586894 108854 622338
rect 108234 586658 108266 586894
rect 108502 586658 108586 586894
rect 108822 586658 108854 586894
rect 108234 586574 108854 586658
rect 108234 586338 108266 586574
rect 108502 586338 108586 586574
rect 108822 586338 108854 586574
rect 108234 550894 108854 586338
rect 108234 550658 108266 550894
rect 108502 550658 108586 550894
rect 108822 550658 108854 550894
rect 108234 550574 108854 550658
rect 108234 550338 108266 550574
rect 108502 550338 108586 550574
rect 108822 550338 108854 550574
rect 108234 514894 108854 550338
rect 108234 514658 108266 514894
rect 108502 514658 108586 514894
rect 108822 514658 108854 514894
rect 108234 514574 108854 514658
rect 108234 514338 108266 514574
rect 108502 514338 108586 514574
rect 108822 514338 108854 514574
rect 108234 478894 108854 514338
rect 108234 478658 108266 478894
rect 108502 478658 108586 478894
rect 108822 478658 108854 478894
rect 108234 478574 108854 478658
rect 108234 478338 108266 478574
rect 108502 478338 108586 478574
rect 108822 478338 108854 478574
rect 108234 442894 108854 478338
rect 108234 442658 108266 442894
rect 108502 442658 108586 442894
rect 108822 442658 108854 442894
rect 108234 442574 108854 442658
rect 108234 442338 108266 442574
rect 108502 442338 108586 442574
rect 108822 442338 108854 442574
rect 108234 406894 108854 442338
rect 108234 406658 108266 406894
rect 108502 406658 108586 406894
rect 108822 406658 108854 406894
rect 108234 406574 108854 406658
rect 108234 406338 108266 406574
rect 108502 406338 108586 406574
rect 108822 406338 108854 406574
rect 108234 370894 108854 406338
rect 108234 370658 108266 370894
rect 108502 370658 108586 370894
rect 108822 370658 108854 370894
rect 108234 370574 108854 370658
rect 108234 370338 108266 370574
rect 108502 370338 108586 370574
rect 108822 370338 108854 370574
rect 108234 334894 108854 370338
rect 108234 334658 108266 334894
rect 108502 334658 108586 334894
rect 108822 334658 108854 334894
rect 108234 334574 108854 334658
rect 108234 334338 108266 334574
rect 108502 334338 108586 334574
rect 108822 334338 108854 334574
rect 108234 298894 108854 334338
rect 108234 298658 108266 298894
rect 108502 298658 108586 298894
rect 108822 298658 108854 298894
rect 108234 298574 108854 298658
rect 108234 298338 108266 298574
rect 108502 298338 108586 298574
rect 108822 298338 108854 298574
rect 108234 262894 108854 298338
rect 108234 262658 108266 262894
rect 108502 262658 108586 262894
rect 108822 262658 108854 262894
rect 108234 262574 108854 262658
rect 108234 262338 108266 262574
rect 108502 262338 108586 262574
rect 108822 262338 108854 262574
rect 108234 226894 108854 262338
rect 108234 226658 108266 226894
rect 108502 226658 108586 226894
rect 108822 226658 108854 226894
rect 108234 226574 108854 226658
rect 108234 226338 108266 226574
rect 108502 226338 108586 226574
rect 108822 226338 108854 226574
rect 108234 190894 108854 226338
rect 108234 190658 108266 190894
rect 108502 190658 108586 190894
rect 108822 190658 108854 190894
rect 108234 190574 108854 190658
rect 108234 190338 108266 190574
rect 108502 190338 108586 190574
rect 108822 190338 108854 190574
rect 108234 154894 108854 190338
rect 108234 154658 108266 154894
rect 108502 154658 108586 154894
rect 108822 154658 108854 154894
rect 108234 154574 108854 154658
rect 108234 154338 108266 154574
rect 108502 154338 108586 154574
rect 108822 154338 108854 154574
rect 108234 118894 108854 154338
rect 108234 118658 108266 118894
rect 108502 118658 108586 118894
rect 108822 118658 108854 118894
rect 108234 118574 108854 118658
rect 108234 118338 108266 118574
rect 108502 118338 108586 118574
rect 108822 118338 108854 118574
rect 108234 82894 108854 118338
rect 108234 82658 108266 82894
rect 108502 82658 108586 82894
rect 108822 82658 108854 82894
rect 108234 82574 108854 82658
rect 108234 82338 108266 82574
rect 108502 82338 108586 82574
rect 108822 82338 108854 82574
rect 108234 46894 108854 82338
rect 108234 46658 108266 46894
rect 108502 46658 108586 46894
rect 108822 46658 108854 46894
rect 108234 46574 108854 46658
rect 108234 46338 108266 46574
rect 108502 46338 108586 46574
rect 108822 46338 108854 46574
rect 108234 10894 108854 46338
rect 108234 10658 108266 10894
rect 108502 10658 108586 10894
rect 108822 10658 108854 10894
rect 108234 10574 108854 10658
rect 108234 10338 108266 10574
rect 108502 10338 108586 10574
rect 108822 10338 108854 10574
rect 108234 -4186 108854 10338
rect 110794 705798 111414 705830
rect 110794 705562 110826 705798
rect 111062 705562 111146 705798
rect 111382 705562 111414 705798
rect 110794 705478 111414 705562
rect 110794 705242 110826 705478
rect 111062 705242 111146 705478
rect 111382 705242 111414 705478
rect 110794 669454 111414 705242
rect 110794 669218 110826 669454
rect 111062 669218 111146 669454
rect 111382 669218 111414 669454
rect 110794 669134 111414 669218
rect 110794 668898 110826 669134
rect 111062 668898 111146 669134
rect 111382 668898 111414 669134
rect 110794 633454 111414 668898
rect 110794 633218 110826 633454
rect 111062 633218 111146 633454
rect 111382 633218 111414 633454
rect 110794 633134 111414 633218
rect 110794 632898 110826 633134
rect 111062 632898 111146 633134
rect 111382 632898 111414 633134
rect 110794 597454 111414 632898
rect 110794 597218 110826 597454
rect 111062 597218 111146 597454
rect 111382 597218 111414 597454
rect 110794 597134 111414 597218
rect 110794 596898 110826 597134
rect 111062 596898 111146 597134
rect 111382 596898 111414 597134
rect 110794 561454 111414 596898
rect 110794 561218 110826 561454
rect 111062 561218 111146 561454
rect 111382 561218 111414 561454
rect 110794 561134 111414 561218
rect 110794 560898 110826 561134
rect 111062 560898 111146 561134
rect 111382 560898 111414 561134
rect 110794 525454 111414 560898
rect 110794 525218 110826 525454
rect 111062 525218 111146 525454
rect 111382 525218 111414 525454
rect 110794 525134 111414 525218
rect 110794 524898 110826 525134
rect 111062 524898 111146 525134
rect 111382 524898 111414 525134
rect 110794 489454 111414 524898
rect 110794 489218 110826 489454
rect 111062 489218 111146 489454
rect 111382 489218 111414 489454
rect 110794 489134 111414 489218
rect 110794 488898 110826 489134
rect 111062 488898 111146 489134
rect 111382 488898 111414 489134
rect 110794 453454 111414 488898
rect 110794 453218 110826 453454
rect 111062 453218 111146 453454
rect 111382 453218 111414 453454
rect 110794 453134 111414 453218
rect 110794 452898 110826 453134
rect 111062 452898 111146 453134
rect 111382 452898 111414 453134
rect 110794 417454 111414 452898
rect 110794 417218 110826 417454
rect 111062 417218 111146 417454
rect 111382 417218 111414 417454
rect 110794 417134 111414 417218
rect 110794 416898 110826 417134
rect 111062 416898 111146 417134
rect 111382 416898 111414 417134
rect 110794 381454 111414 416898
rect 110794 381218 110826 381454
rect 111062 381218 111146 381454
rect 111382 381218 111414 381454
rect 110794 381134 111414 381218
rect 110794 380898 110826 381134
rect 111062 380898 111146 381134
rect 111382 380898 111414 381134
rect 110794 345454 111414 380898
rect 110794 345218 110826 345454
rect 111062 345218 111146 345454
rect 111382 345218 111414 345454
rect 110794 345134 111414 345218
rect 110794 344898 110826 345134
rect 111062 344898 111146 345134
rect 111382 344898 111414 345134
rect 110794 309454 111414 344898
rect 110794 309218 110826 309454
rect 111062 309218 111146 309454
rect 111382 309218 111414 309454
rect 110794 309134 111414 309218
rect 110794 308898 110826 309134
rect 111062 308898 111146 309134
rect 111382 308898 111414 309134
rect 110794 273454 111414 308898
rect 110794 273218 110826 273454
rect 111062 273218 111146 273454
rect 111382 273218 111414 273454
rect 110794 273134 111414 273218
rect 110794 272898 110826 273134
rect 111062 272898 111146 273134
rect 111382 272898 111414 273134
rect 110794 237454 111414 272898
rect 110794 237218 110826 237454
rect 111062 237218 111146 237454
rect 111382 237218 111414 237454
rect 110794 237134 111414 237218
rect 110794 236898 110826 237134
rect 111062 236898 111146 237134
rect 111382 236898 111414 237134
rect 110794 201454 111414 236898
rect 110794 201218 110826 201454
rect 111062 201218 111146 201454
rect 111382 201218 111414 201454
rect 110794 201134 111414 201218
rect 110794 200898 110826 201134
rect 111062 200898 111146 201134
rect 111382 200898 111414 201134
rect 110794 165454 111414 200898
rect 110794 165218 110826 165454
rect 111062 165218 111146 165454
rect 111382 165218 111414 165454
rect 110794 165134 111414 165218
rect 110794 164898 110826 165134
rect 111062 164898 111146 165134
rect 111382 164898 111414 165134
rect 110794 129454 111414 164898
rect 110794 129218 110826 129454
rect 111062 129218 111146 129454
rect 111382 129218 111414 129454
rect 110794 129134 111414 129218
rect 110794 128898 110826 129134
rect 111062 128898 111146 129134
rect 111382 128898 111414 129134
rect 110794 93454 111414 128898
rect 110794 93218 110826 93454
rect 111062 93218 111146 93454
rect 111382 93218 111414 93454
rect 110794 93134 111414 93218
rect 110794 92898 110826 93134
rect 111062 92898 111146 93134
rect 111382 92898 111414 93134
rect 110794 57454 111414 92898
rect 110794 57218 110826 57454
rect 111062 57218 111146 57454
rect 111382 57218 111414 57454
rect 110794 57134 111414 57218
rect 110794 56898 110826 57134
rect 111062 56898 111146 57134
rect 111382 56898 111414 57134
rect 110794 21454 111414 56898
rect 110794 21218 110826 21454
rect 111062 21218 111146 21454
rect 111382 21218 111414 21454
rect 110794 21134 111414 21218
rect 110794 20898 110826 21134
rect 111062 20898 111146 21134
rect 111382 20898 111414 21134
rect 110794 -1306 111414 20898
rect 110794 -1542 110826 -1306
rect 111062 -1542 111146 -1306
rect 111382 -1542 111414 -1306
rect 110794 -1626 111414 -1542
rect 110794 -1862 110826 -1626
rect 111062 -1862 111146 -1626
rect 111382 -1862 111414 -1626
rect 110794 -1894 111414 -1862
rect 111954 698614 112574 710042
rect 121954 711558 122574 711590
rect 121954 711322 121986 711558
rect 122222 711322 122306 711558
rect 122542 711322 122574 711558
rect 121954 711238 122574 711322
rect 121954 711002 121986 711238
rect 122222 711002 122306 711238
rect 122542 711002 122574 711238
rect 118234 709638 118854 709670
rect 118234 709402 118266 709638
rect 118502 709402 118586 709638
rect 118822 709402 118854 709638
rect 118234 709318 118854 709402
rect 118234 709082 118266 709318
rect 118502 709082 118586 709318
rect 118822 709082 118854 709318
rect 111954 698378 111986 698614
rect 112222 698378 112306 698614
rect 112542 698378 112574 698614
rect 111954 698294 112574 698378
rect 111954 698058 111986 698294
rect 112222 698058 112306 698294
rect 112542 698058 112574 698294
rect 111954 662614 112574 698058
rect 111954 662378 111986 662614
rect 112222 662378 112306 662614
rect 112542 662378 112574 662614
rect 111954 662294 112574 662378
rect 111954 662058 111986 662294
rect 112222 662058 112306 662294
rect 112542 662058 112574 662294
rect 111954 626614 112574 662058
rect 111954 626378 111986 626614
rect 112222 626378 112306 626614
rect 112542 626378 112574 626614
rect 111954 626294 112574 626378
rect 111954 626058 111986 626294
rect 112222 626058 112306 626294
rect 112542 626058 112574 626294
rect 111954 590614 112574 626058
rect 111954 590378 111986 590614
rect 112222 590378 112306 590614
rect 112542 590378 112574 590614
rect 111954 590294 112574 590378
rect 111954 590058 111986 590294
rect 112222 590058 112306 590294
rect 112542 590058 112574 590294
rect 111954 554614 112574 590058
rect 111954 554378 111986 554614
rect 112222 554378 112306 554614
rect 112542 554378 112574 554614
rect 111954 554294 112574 554378
rect 111954 554058 111986 554294
rect 112222 554058 112306 554294
rect 112542 554058 112574 554294
rect 111954 518614 112574 554058
rect 111954 518378 111986 518614
rect 112222 518378 112306 518614
rect 112542 518378 112574 518614
rect 111954 518294 112574 518378
rect 111954 518058 111986 518294
rect 112222 518058 112306 518294
rect 112542 518058 112574 518294
rect 111954 482614 112574 518058
rect 111954 482378 111986 482614
rect 112222 482378 112306 482614
rect 112542 482378 112574 482614
rect 111954 482294 112574 482378
rect 111954 482058 111986 482294
rect 112222 482058 112306 482294
rect 112542 482058 112574 482294
rect 111954 446614 112574 482058
rect 111954 446378 111986 446614
rect 112222 446378 112306 446614
rect 112542 446378 112574 446614
rect 111954 446294 112574 446378
rect 111954 446058 111986 446294
rect 112222 446058 112306 446294
rect 112542 446058 112574 446294
rect 111954 410614 112574 446058
rect 111954 410378 111986 410614
rect 112222 410378 112306 410614
rect 112542 410378 112574 410614
rect 111954 410294 112574 410378
rect 111954 410058 111986 410294
rect 112222 410058 112306 410294
rect 112542 410058 112574 410294
rect 111954 374614 112574 410058
rect 111954 374378 111986 374614
rect 112222 374378 112306 374614
rect 112542 374378 112574 374614
rect 111954 374294 112574 374378
rect 111954 374058 111986 374294
rect 112222 374058 112306 374294
rect 112542 374058 112574 374294
rect 111954 338614 112574 374058
rect 111954 338378 111986 338614
rect 112222 338378 112306 338614
rect 112542 338378 112574 338614
rect 111954 338294 112574 338378
rect 111954 338058 111986 338294
rect 112222 338058 112306 338294
rect 112542 338058 112574 338294
rect 111954 302614 112574 338058
rect 111954 302378 111986 302614
rect 112222 302378 112306 302614
rect 112542 302378 112574 302614
rect 111954 302294 112574 302378
rect 111954 302058 111986 302294
rect 112222 302058 112306 302294
rect 112542 302058 112574 302294
rect 111954 266614 112574 302058
rect 111954 266378 111986 266614
rect 112222 266378 112306 266614
rect 112542 266378 112574 266614
rect 111954 266294 112574 266378
rect 111954 266058 111986 266294
rect 112222 266058 112306 266294
rect 112542 266058 112574 266294
rect 111954 230614 112574 266058
rect 111954 230378 111986 230614
rect 112222 230378 112306 230614
rect 112542 230378 112574 230614
rect 111954 230294 112574 230378
rect 111954 230058 111986 230294
rect 112222 230058 112306 230294
rect 112542 230058 112574 230294
rect 111954 194614 112574 230058
rect 111954 194378 111986 194614
rect 112222 194378 112306 194614
rect 112542 194378 112574 194614
rect 111954 194294 112574 194378
rect 111954 194058 111986 194294
rect 112222 194058 112306 194294
rect 112542 194058 112574 194294
rect 111954 158614 112574 194058
rect 111954 158378 111986 158614
rect 112222 158378 112306 158614
rect 112542 158378 112574 158614
rect 111954 158294 112574 158378
rect 111954 158058 111986 158294
rect 112222 158058 112306 158294
rect 112542 158058 112574 158294
rect 111954 122614 112574 158058
rect 111954 122378 111986 122614
rect 112222 122378 112306 122614
rect 112542 122378 112574 122614
rect 111954 122294 112574 122378
rect 111954 122058 111986 122294
rect 112222 122058 112306 122294
rect 112542 122058 112574 122294
rect 111954 86614 112574 122058
rect 111954 86378 111986 86614
rect 112222 86378 112306 86614
rect 112542 86378 112574 86614
rect 111954 86294 112574 86378
rect 111954 86058 111986 86294
rect 112222 86058 112306 86294
rect 112542 86058 112574 86294
rect 111954 50614 112574 86058
rect 111954 50378 111986 50614
rect 112222 50378 112306 50614
rect 112542 50378 112574 50614
rect 111954 50294 112574 50378
rect 111954 50058 111986 50294
rect 112222 50058 112306 50294
rect 112542 50058 112574 50294
rect 111954 14614 112574 50058
rect 111954 14378 111986 14614
rect 112222 14378 112306 14614
rect 112542 14378 112574 14614
rect 111954 14294 112574 14378
rect 111954 14058 111986 14294
rect 112222 14058 112306 14294
rect 112542 14058 112574 14294
rect 108234 -4422 108266 -4186
rect 108502 -4422 108586 -4186
rect 108822 -4422 108854 -4186
rect 108234 -4506 108854 -4422
rect 108234 -4742 108266 -4506
rect 108502 -4742 108586 -4506
rect 108822 -4742 108854 -4506
rect 108234 -5734 108854 -4742
rect 101954 -7302 101986 -7066
rect 102222 -7302 102306 -7066
rect 102542 -7302 102574 -7066
rect 101954 -7386 102574 -7302
rect 101954 -7622 101986 -7386
rect 102222 -7622 102306 -7386
rect 102542 -7622 102574 -7386
rect 101954 -7654 102574 -7622
rect 111954 -6106 112574 14058
rect 114514 707718 115134 707750
rect 114514 707482 114546 707718
rect 114782 707482 114866 707718
rect 115102 707482 115134 707718
rect 114514 707398 115134 707482
rect 114514 707162 114546 707398
rect 114782 707162 114866 707398
rect 115102 707162 115134 707398
rect 114514 673174 115134 707162
rect 114514 672938 114546 673174
rect 114782 672938 114866 673174
rect 115102 672938 115134 673174
rect 114514 672854 115134 672938
rect 114514 672618 114546 672854
rect 114782 672618 114866 672854
rect 115102 672618 115134 672854
rect 114514 637174 115134 672618
rect 114514 636938 114546 637174
rect 114782 636938 114866 637174
rect 115102 636938 115134 637174
rect 114514 636854 115134 636938
rect 114514 636618 114546 636854
rect 114782 636618 114866 636854
rect 115102 636618 115134 636854
rect 114514 601174 115134 636618
rect 114514 600938 114546 601174
rect 114782 600938 114866 601174
rect 115102 600938 115134 601174
rect 114514 600854 115134 600938
rect 114514 600618 114546 600854
rect 114782 600618 114866 600854
rect 115102 600618 115134 600854
rect 114514 565174 115134 600618
rect 114514 564938 114546 565174
rect 114782 564938 114866 565174
rect 115102 564938 115134 565174
rect 114514 564854 115134 564938
rect 114514 564618 114546 564854
rect 114782 564618 114866 564854
rect 115102 564618 115134 564854
rect 114514 529174 115134 564618
rect 114514 528938 114546 529174
rect 114782 528938 114866 529174
rect 115102 528938 115134 529174
rect 114514 528854 115134 528938
rect 114514 528618 114546 528854
rect 114782 528618 114866 528854
rect 115102 528618 115134 528854
rect 114514 493174 115134 528618
rect 114514 492938 114546 493174
rect 114782 492938 114866 493174
rect 115102 492938 115134 493174
rect 114514 492854 115134 492938
rect 114514 492618 114546 492854
rect 114782 492618 114866 492854
rect 115102 492618 115134 492854
rect 114514 457174 115134 492618
rect 114514 456938 114546 457174
rect 114782 456938 114866 457174
rect 115102 456938 115134 457174
rect 114514 456854 115134 456938
rect 114514 456618 114546 456854
rect 114782 456618 114866 456854
rect 115102 456618 115134 456854
rect 114514 421174 115134 456618
rect 114514 420938 114546 421174
rect 114782 420938 114866 421174
rect 115102 420938 115134 421174
rect 114514 420854 115134 420938
rect 114514 420618 114546 420854
rect 114782 420618 114866 420854
rect 115102 420618 115134 420854
rect 114514 385174 115134 420618
rect 114514 384938 114546 385174
rect 114782 384938 114866 385174
rect 115102 384938 115134 385174
rect 114514 384854 115134 384938
rect 114514 384618 114546 384854
rect 114782 384618 114866 384854
rect 115102 384618 115134 384854
rect 114514 349174 115134 384618
rect 114514 348938 114546 349174
rect 114782 348938 114866 349174
rect 115102 348938 115134 349174
rect 114514 348854 115134 348938
rect 114514 348618 114546 348854
rect 114782 348618 114866 348854
rect 115102 348618 115134 348854
rect 114514 313174 115134 348618
rect 114514 312938 114546 313174
rect 114782 312938 114866 313174
rect 115102 312938 115134 313174
rect 114514 312854 115134 312938
rect 114514 312618 114546 312854
rect 114782 312618 114866 312854
rect 115102 312618 115134 312854
rect 114514 277174 115134 312618
rect 114514 276938 114546 277174
rect 114782 276938 114866 277174
rect 115102 276938 115134 277174
rect 114514 276854 115134 276938
rect 114514 276618 114546 276854
rect 114782 276618 114866 276854
rect 115102 276618 115134 276854
rect 114514 241174 115134 276618
rect 114514 240938 114546 241174
rect 114782 240938 114866 241174
rect 115102 240938 115134 241174
rect 114514 240854 115134 240938
rect 114514 240618 114546 240854
rect 114782 240618 114866 240854
rect 115102 240618 115134 240854
rect 114514 205174 115134 240618
rect 114514 204938 114546 205174
rect 114782 204938 114866 205174
rect 115102 204938 115134 205174
rect 114514 204854 115134 204938
rect 114514 204618 114546 204854
rect 114782 204618 114866 204854
rect 115102 204618 115134 204854
rect 114514 169174 115134 204618
rect 114514 168938 114546 169174
rect 114782 168938 114866 169174
rect 115102 168938 115134 169174
rect 114514 168854 115134 168938
rect 114514 168618 114546 168854
rect 114782 168618 114866 168854
rect 115102 168618 115134 168854
rect 114514 133174 115134 168618
rect 114514 132938 114546 133174
rect 114782 132938 114866 133174
rect 115102 132938 115134 133174
rect 114514 132854 115134 132938
rect 114514 132618 114546 132854
rect 114782 132618 114866 132854
rect 115102 132618 115134 132854
rect 114514 97174 115134 132618
rect 114514 96938 114546 97174
rect 114782 96938 114866 97174
rect 115102 96938 115134 97174
rect 114514 96854 115134 96938
rect 114514 96618 114546 96854
rect 114782 96618 114866 96854
rect 115102 96618 115134 96854
rect 114514 61174 115134 96618
rect 114514 60938 114546 61174
rect 114782 60938 114866 61174
rect 115102 60938 115134 61174
rect 114514 60854 115134 60938
rect 114514 60618 114546 60854
rect 114782 60618 114866 60854
rect 115102 60618 115134 60854
rect 114514 25174 115134 60618
rect 114514 24938 114546 25174
rect 114782 24938 114866 25174
rect 115102 24938 115134 25174
rect 114514 24854 115134 24938
rect 114514 24618 114546 24854
rect 114782 24618 114866 24854
rect 115102 24618 115134 24854
rect 114514 -3226 115134 24618
rect 114514 -3462 114546 -3226
rect 114782 -3462 114866 -3226
rect 115102 -3462 115134 -3226
rect 114514 -3546 115134 -3462
rect 114514 -3782 114546 -3546
rect 114782 -3782 114866 -3546
rect 115102 -3782 115134 -3546
rect 114514 -3814 115134 -3782
rect 118234 676894 118854 709082
rect 118234 676658 118266 676894
rect 118502 676658 118586 676894
rect 118822 676658 118854 676894
rect 118234 676574 118854 676658
rect 118234 676338 118266 676574
rect 118502 676338 118586 676574
rect 118822 676338 118854 676574
rect 118234 640894 118854 676338
rect 118234 640658 118266 640894
rect 118502 640658 118586 640894
rect 118822 640658 118854 640894
rect 118234 640574 118854 640658
rect 118234 640338 118266 640574
rect 118502 640338 118586 640574
rect 118822 640338 118854 640574
rect 118234 604894 118854 640338
rect 118234 604658 118266 604894
rect 118502 604658 118586 604894
rect 118822 604658 118854 604894
rect 118234 604574 118854 604658
rect 118234 604338 118266 604574
rect 118502 604338 118586 604574
rect 118822 604338 118854 604574
rect 118234 568894 118854 604338
rect 118234 568658 118266 568894
rect 118502 568658 118586 568894
rect 118822 568658 118854 568894
rect 118234 568574 118854 568658
rect 118234 568338 118266 568574
rect 118502 568338 118586 568574
rect 118822 568338 118854 568574
rect 118234 532894 118854 568338
rect 118234 532658 118266 532894
rect 118502 532658 118586 532894
rect 118822 532658 118854 532894
rect 118234 532574 118854 532658
rect 118234 532338 118266 532574
rect 118502 532338 118586 532574
rect 118822 532338 118854 532574
rect 118234 496894 118854 532338
rect 118234 496658 118266 496894
rect 118502 496658 118586 496894
rect 118822 496658 118854 496894
rect 118234 496574 118854 496658
rect 118234 496338 118266 496574
rect 118502 496338 118586 496574
rect 118822 496338 118854 496574
rect 118234 460894 118854 496338
rect 118234 460658 118266 460894
rect 118502 460658 118586 460894
rect 118822 460658 118854 460894
rect 118234 460574 118854 460658
rect 118234 460338 118266 460574
rect 118502 460338 118586 460574
rect 118822 460338 118854 460574
rect 118234 424894 118854 460338
rect 118234 424658 118266 424894
rect 118502 424658 118586 424894
rect 118822 424658 118854 424894
rect 118234 424574 118854 424658
rect 118234 424338 118266 424574
rect 118502 424338 118586 424574
rect 118822 424338 118854 424574
rect 118234 388894 118854 424338
rect 118234 388658 118266 388894
rect 118502 388658 118586 388894
rect 118822 388658 118854 388894
rect 118234 388574 118854 388658
rect 118234 388338 118266 388574
rect 118502 388338 118586 388574
rect 118822 388338 118854 388574
rect 118234 352894 118854 388338
rect 118234 352658 118266 352894
rect 118502 352658 118586 352894
rect 118822 352658 118854 352894
rect 118234 352574 118854 352658
rect 118234 352338 118266 352574
rect 118502 352338 118586 352574
rect 118822 352338 118854 352574
rect 118234 316894 118854 352338
rect 118234 316658 118266 316894
rect 118502 316658 118586 316894
rect 118822 316658 118854 316894
rect 118234 316574 118854 316658
rect 118234 316338 118266 316574
rect 118502 316338 118586 316574
rect 118822 316338 118854 316574
rect 118234 280894 118854 316338
rect 118234 280658 118266 280894
rect 118502 280658 118586 280894
rect 118822 280658 118854 280894
rect 118234 280574 118854 280658
rect 118234 280338 118266 280574
rect 118502 280338 118586 280574
rect 118822 280338 118854 280574
rect 118234 244894 118854 280338
rect 118234 244658 118266 244894
rect 118502 244658 118586 244894
rect 118822 244658 118854 244894
rect 118234 244574 118854 244658
rect 118234 244338 118266 244574
rect 118502 244338 118586 244574
rect 118822 244338 118854 244574
rect 118234 208894 118854 244338
rect 118234 208658 118266 208894
rect 118502 208658 118586 208894
rect 118822 208658 118854 208894
rect 118234 208574 118854 208658
rect 118234 208338 118266 208574
rect 118502 208338 118586 208574
rect 118822 208338 118854 208574
rect 118234 172894 118854 208338
rect 118234 172658 118266 172894
rect 118502 172658 118586 172894
rect 118822 172658 118854 172894
rect 118234 172574 118854 172658
rect 118234 172338 118266 172574
rect 118502 172338 118586 172574
rect 118822 172338 118854 172574
rect 118234 136894 118854 172338
rect 118234 136658 118266 136894
rect 118502 136658 118586 136894
rect 118822 136658 118854 136894
rect 118234 136574 118854 136658
rect 118234 136338 118266 136574
rect 118502 136338 118586 136574
rect 118822 136338 118854 136574
rect 118234 100894 118854 136338
rect 118234 100658 118266 100894
rect 118502 100658 118586 100894
rect 118822 100658 118854 100894
rect 118234 100574 118854 100658
rect 118234 100338 118266 100574
rect 118502 100338 118586 100574
rect 118822 100338 118854 100574
rect 118234 64894 118854 100338
rect 118234 64658 118266 64894
rect 118502 64658 118586 64894
rect 118822 64658 118854 64894
rect 118234 64574 118854 64658
rect 118234 64338 118266 64574
rect 118502 64338 118586 64574
rect 118822 64338 118854 64574
rect 118234 28894 118854 64338
rect 118234 28658 118266 28894
rect 118502 28658 118586 28894
rect 118822 28658 118854 28894
rect 118234 28574 118854 28658
rect 118234 28338 118266 28574
rect 118502 28338 118586 28574
rect 118822 28338 118854 28574
rect 118234 -5146 118854 28338
rect 120794 704838 121414 705830
rect 120794 704602 120826 704838
rect 121062 704602 121146 704838
rect 121382 704602 121414 704838
rect 120794 704518 121414 704602
rect 120794 704282 120826 704518
rect 121062 704282 121146 704518
rect 121382 704282 121414 704518
rect 120794 687454 121414 704282
rect 120794 687218 120826 687454
rect 121062 687218 121146 687454
rect 121382 687218 121414 687454
rect 120794 687134 121414 687218
rect 120794 686898 120826 687134
rect 121062 686898 121146 687134
rect 121382 686898 121414 687134
rect 120794 651454 121414 686898
rect 120794 651218 120826 651454
rect 121062 651218 121146 651454
rect 121382 651218 121414 651454
rect 120794 651134 121414 651218
rect 120794 650898 120826 651134
rect 121062 650898 121146 651134
rect 121382 650898 121414 651134
rect 120794 615454 121414 650898
rect 120794 615218 120826 615454
rect 121062 615218 121146 615454
rect 121382 615218 121414 615454
rect 120794 615134 121414 615218
rect 120794 614898 120826 615134
rect 121062 614898 121146 615134
rect 121382 614898 121414 615134
rect 120794 579454 121414 614898
rect 120794 579218 120826 579454
rect 121062 579218 121146 579454
rect 121382 579218 121414 579454
rect 120794 579134 121414 579218
rect 120794 578898 120826 579134
rect 121062 578898 121146 579134
rect 121382 578898 121414 579134
rect 120794 543454 121414 578898
rect 120794 543218 120826 543454
rect 121062 543218 121146 543454
rect 121382 543218 121414 543454
rect 120794 543134 121414 543218
rect 120794 542898 120826 543134
rect 121062 542898 121146 543134
rect 121382 542898 121414 543134
rect 120794 507454 121414 542898
rect 120794 507218 120826 507454
rect 121062 507218 121146 507454
rect 121382 507218 121414 507454
rect 120794 507134 121414 507218
rect 120794 506898 120826 507134
rect 121062 506898 121146 507134
rect 121382 506898 121414 507134
rect 120794 471454 121414 506898
rect 120794 471218 120826 471454
rect 121062 471218 121146 471454
rect 121382 471218 121414 471454
rect 120794 471134 121414 471218
rect 120794 470898 120826 471134
rect 121062 470898 121146 471134
rect 121382 470898 121414 471134
rect 120794 435454 121414 470898
rect 120794 435218 120826 435454
rect 121062 435218 121146 435454
rect 121382 435218 121414 435454
rect 120794 435134 121414 435218
rect 120794 434898 120826 435134
rect 121062 434898 121146 435134
rect 121382 434898 121414 435134
rect 120794 399454 121414 434898
rect 120794 399218 120826 399454
rect 121062 399218 121146 399454
rect 121382 399218 121414 399454
rect 120794 399134 121414 399218
rect 120794 398898 120826 399134
rect 121062 398898 121146 399134
rect 121382 398898 121414 399134
rect 120794 363454 121414 398898
rect 120794 363218 120826 363454
rect 121062 363218 121146 363454
rect 121382 363218 121414 363454
rect 120794 363134 121414 363218
rect 120794 362898 120826 363134
rect 121062 362898 121146 363134
rect 121382 362898 121414 363134
rect 120794 327454 121414 362898
rect 120794 327218 120826 327454
rect 121062 327218 121146 327454
rect 121382 327218 121414 327454
rect 120794 327134 121414 327218
rect 120794 326898 120826 327134
rect 121062 326898 121146 327134
rect 121382 326898 121414 327134
rect 120794 291454 121414 326898
rect 120794 291218 120826 291454
rect 121062 291218 121146 291454
rect 121382 291218 121414 291454
rect 120794 291134 121414 291218
rect 120794 290898 120826 291134
rect 121062 290898 121146 291134
rect 121382 290898 121414 291134
rect 120794 255454 121414 290898
rect 120794 255218 120826 255454
rect 121062 255218 121146 255454
rect 121382 255218 121414 255454
rect 120794 255134 121414 255218
rect 120794 254898 120826 255134
rect 121062 254898 121146 255134
rect 121382 254898 121414 255134
rect 120794 219454 121414 254898
rect 120794 219218 120826 219454
rect 121062 219218 121146 219454
rect 121382 219218 121414 219454
rect 120794 219134 121414 219218
rect 120794 218898 120826 219134
rect 121062 218898 121146 219134
rect 121382 218898 121414 219134
rect 120794 183454 121414 218898
rect 120794 183218 120826 183454
rect 121062 183218 121146 183454
rect 121382 183218 121414 183454
rect 120794 183134 121414 183218
rect 120794 182898 120826 183134
rect 121062 182898 121146 183134
rect 121382 182898 121414 183134
rect 120794 147454 121414 182898
rect 120794 147218 120826 147454
rect 121062 147218 121146 147454
rect 121382 147218 121414 147454
rect 120794 147134 121414 147218
rect 120794 146898 120826 147134
rect 121062 146898 121146 147134
rect 121382 146898 121414 147134
rect 120794 111454 121414 146898
rect 120794 111218 120826 111454
rect 121062 111218 121146 111454
rect 121382 111218 121414 111454
rect 120794 111134 121414 111218
rect 120794 110898 120826 111134
rect 121062 110898 121146 111134
rect 121382 110898 121414 111134
rect 120794 75454 121414 110898
rect 120794 75218 120826 75454
rect 121062 75218 121146 75454
rect 121382 75218 121414 75454
rect 120794 75134 121414 75218
rect 120794 74898 120826 75134
rect 121062 74898 121146 75134
rect 121382 74898 121414 75134
rect 120794 39454 121414 74898
rect 120794 39218 120826 39454
rect 121062 39218 121146 39454
rect 121382 39218 121414 39454
rect 120794 39134 121414 39218
rect 120794 38898 120826 39134
rect 121062 38898 121146 39134
rect 121382 38898 121414 39134
rect 120794 3454 121414 38898
rect 120794 3218 120826 3454
rect 121062 3218 121146 3454
rect 121382 3218 121414 3454
rect 120794 3134 121414 3218
rect 120794 2898 120826 3134
rect 121062 2898 121146 3134
rect 121382 2898 121414 3134
rect 120794 -346 121414 2898
rect 120794 -582 120826 -346
rect 121062 -582 121146 -346
rect 121382 -582 121414 -346
rect 120794 -666 121414 -582
rect 120794 -902 120826 -666
rect 121062 -902 121146 -666
rect 121382 -902 121414 -666
rect 120794 -1894 121414 -902
rect 121954 680614 122574 711002
rect 131954 710598 132574 711590
rect 131954 710362 131986 710598
rect 132222 710362 132306 710598
rect 132542 710362 132574 710598
rect 131954 710278 132574 710362
rect 131954 710042 131986 710278
rect 132222 710042 132306 710278
rect 132542 710042 132574 710278
rect 128234 708678 128854 709670
rect 128234 708442 128266 708678
rect 128502 708442 128586 708678
rect 128822 708442 128854 708678
rect 128234 708358 128854 708442
rect 128234 708122 128266 708358
rect 128502 708122 128586 708358
rect 128822 708122 128854 708358
rect 121954 680378 121986 680614
rect 122222 680378 122306 680614
rect 122542 680378 122574 680614
rect 121954 680294 122574 680378
rect 121954 680058 121986 680294
rect 122222 680058 122306 680294
rect 122542 680058 122574 680294
rect 121954 644614 122574 680058
rect 121954 644378 121986 644614
rect 122222 644378 122306 644614
rect 122542 644378 122574 644614
rect 121954 644294 122574 644378
rect 121954 644058 121986 644294
rect 122222 644058 122306 644294
rect 122542 644058 122574 644294
rect 121954 608614 122574 644058
rect 121954 608378 121986 608614
rect 122222 608378 122306 608614
rect 122542 608378 122574 608614
rect 121954 608294 122574 608378
rect 121954 608058 121986 608294
rect 122222 608058 122306 608294
rect 122542 608058 122574 608294
rect 121954 572614 122574 608058
rect 121954 572378 121986 572614
rect 122222 572378 122306 572614
rect 122542 572378 122574 572614
rect 121954 572294 122574 572378
rect 121954 572058 121986 572294
rect 122222 572058 122306 572294
rect 122542 572058 122574 572294
rect 121954 536614 122574 572058
rect 121954 536378 121986 536614
rect 122222 536378 122306 536614
rect 122542 536378 122574 536614
rect 121954 536294 122574 536378
rect 121954 536058 121986 536294
rect 122222 536058 122306 536294
rect 122542 536058 122574 536294
rect 121954 500614 122574 536058
rect 121954 500378 121986 500614
rect 122222 500378 122306 500614
rect 122542 500378 122574 500614
rect 121954 500294 122574 500378
rect 121954 500058 121986 500294
rect 122222 500058 122306 500294
rect 122542 500058 122574 500294
rect 121954 464614 122574 500058
rect 121954 464378 121986 464614
rect 122222 464378 122306 464614
rect 122542 464378 122574 464614
rect 121954 464294 122574 464378
rect 121954 464058 121986 464294
rect 122222 464058 122306 464294
rect 122542 464058 122574 464294
rect 121954 428614 122574 464058
rect 121954 428378 121986 428614
rect 122222 428378 122306 428614
rect 122542 428378 122574 428614
rect 121954 428294 122574 428378
rect 121954 428058 121986 428294
rect 122222 428058 122306 428294
rect 122542 428058 122574 428294
rect 121954 392614 122574 428058
rect 121954 392378 121986 392614
rect 122222 392378 122306 392614
rect 122542 392378 122574 392614
rect 121954 392294 122574 392378
rect 121954 392058 121986 392294
rect 122222 392058 122306 392294
rect 122542 392058 122574 392294
rect 121954 356614 122574 392058
rect 121954 356378 121986 356614
rect 122222 356378 122306 356614
rect 122542 356378 122574 356614
rect 121954 356294 122574 356378
rect 121954 356058 121986 356294
rect 122222 356058 122306 356294
rect 122542 356058 122574 356294
rect 121954 320614 122574 356058
rect 121954 320378 121986 320614
rect 122222 320378 122306 320614
rect 122542 320378 122574 320614
rect 121954 320294 122574 320378
rect 121954 320058 121986 320294
rect 122222 320058 122306 320294
rect 122542 320058 122574 320294
rect 121954 284614 122574 320058
rect 121954 284378 121986 284614
rect 122222 284378 122306 284614
rect 122542 284378 122574 284614
rect 121954 284294 122574 284378
rect 121954 284058 121986 284294
rect 122222 284058 122306 284294
rect 122542 284058 122574 284294
rect 121954 248614 122574 284058
rect 121954 248378 121986 248614
rect 122222 248378 122306 248614
rect 122542 248378 122574 248614
rect 121954 248294 122574 248378
rect 121954 248058 121986 248294
rect 122222 248058 122306 248294
rect 122542 248058 122574 248294
rect 121954 212614 122574 248058
rect 121954 212378 121986 212614
rect 122222 212378 122306 212614
rect 122542 212378 122574 212614
rect 121954 212294 122574 212378
rect 121954 212058 121986 212294
rect 122222 212058 122306 212294
rect 122542 212058 122574 212294
rect 121954 176614 122574 212058
rect 121954 176378 121986 176614
rect 122222 176378 122306 176614
rect 122542 176378 122574 176614
rect 121954 176294 122574 176378
rect 121954 176058 121986 176294
rect 122222 176058 122306 176294
rect 122542 176058 122574 176294
rect 121954 140614 122574 176058
rect 121954 140378 121986 140614
rect 122222 140378 122306 140614
rect 122542 140378 122574 140614
rect 121954 140294 122574 140378
rect 121954 140058 121986 140294
rect 122222 140058 122306 140294
rect 122542 140058 122574 140294
rect 121954 104614 122574 140058
rect 121954 104378 121986 104614
rect 122222 104378 122306 104614
rect 122542 104378 122574 104614
rect 121954 104294 122574 104378
rect 121954 104058 121986 104294
rect 122222 104058 122306 104294
rect 122542 104058 122574 104294
rect 121954 68614 122574 104058
rect 121954 68378 121986 68614
rect 122222 68378 122306 68614
rect 122542 68378 122574 68614
rect 121954 68294 122574 68378
rect 121954 68058 121986 68294
rect 122222 68058 122306 68294
rect 122542 68058 122574 68294
rect 121954 32614 122574 68058
rect 121954 32378 121986 32614
rect 122222 32378 122306 32614
rect 122542 32378 122574 32614
rect 121954 32294 122574 32378
rect 121954 32058 121986 32294
rect 122222 32058 122306 32294
rect 122542 32058 122574 32294
rect 118234 -5382 118266 -5146
rect 118502 -5382 118586 -5146
rect 118822 -5382 118854 -5146
rect 118234 -5466 118854 -5382
rect 118234 -5702 118266 -5466
rect 118502 -5702 118586 -5466
rect 118822 -5702 118854 -5466
rect 118234 -5734 118854 -5702
rect 111954 -6342 111986 -6106
rect 112222 -6342 112306 -6106
rect 112542 -6342 112574 -6106
rect 111954 -6426 112574 -6342
rect 111954 -6662 111986 -6426
rect 112222 -6662 112306 -6426
rect 112542 -6662 112574 -6426
rect 111954 -7654 112574 -6662
rect 121954 -7066 122574 32058
rect 124514 706758 125134 707750
rect 124514 706522 124546 706758
rect 124782 706522 124866 706758
rect 125102 706522 125134 706758
rect 124514 706438 125134 706522
rect 124514 706202 124546 706438
rect 124782 706202 124866 706438
rect 125102 706202 125134 706438
rect 124514 691174 125134 706202
rect 124514 690938 124546 691174
rect 124782 690938 124866 691174
rect 125102 690938 125134 691174
rect 124514 690854 125134 690938
rect 124514 690618 124546 690854
rect 124782 690618 124866 690854
rect 125102 690618 125134 690854
rect 124514 655174 125134 690618
rect 124514 654938 124546 655174
rect 124782 654938 124866 655174
rect 125102 654938 125134 655174
rect 124514 654854 125134 654938
rect 124514 654618 124546 654854
rect 124782 654618 124866 654854
rect 125102 654618 125134 654854
rect 124514 619174 125134 654618
rect 124514 618938 124546 619174
rect 124782 618938 124866 619174
rect 125102 618938 125134 619174
rect 124514 618854 125134 618938
rect 124514 618618 124546 618854
rect 124782 618618 124866 618854
rect 125102 618618 125134 618854
rect 124514 583174 125134 618618
rect 124514 582938 124546 583174
rect 124782 582938 124866 583174
rect 125102 582938 125134 583174
rect 124514 582854 125134 582938
rect 124514 582618 124546 582854
rect 124782 582618 124866 582854
rect 125102 582618 125134 582854
rect 124514 547174 125134 582618
rect 124514 546938 124546 547174
rect 124782 546938 124866 547174
rect 125102 546938 125134 547174
rect 124514 546854 125134 546938
rect 124514 546618 124546 546854
rect 124782 546618 124866 546854
rect 125102 546618 125134 546854
rect 124514 511174 125134 546618
rect 124514 510938 124546 511174
rect 124782 510938 124866 511174
rect 125102 510938 125134 511174
rect 124514 510854 125134 510938
rect 124514 510618 124546 510854
rect 124782 510618 124866 510854
rect 125102 510618 125134 510854
rect 124514 475174 125134 510618
rect 124514 474938 124546 475174
rect 124782 474938 124866 475174
rect 125102 474938 125134 475174
rect 124514 474854 125134 474938
rect 124514 474618 124546 474854
rect 124782 474618 124866 474854
rect 125102 474618 125134 474854
rect 124514 439174 125134 474618
rect 124514 438938 124546 439174
rect 124782 438938 124866 439174
rect 125102 438938 125134 439174
rect 124514 438854 125134 438938
rect 124514 438618 124546 438854
rect 124782 438618 124866 438854
rect 125102 438618 125134 438854
rect 124514 403174 125134 438618
rect 124514 402938 124546 403174
rect 124782 402938 124866 403174
rect 125102 402938 125134 403174
rect 124514 402854 125134 402938
rect 124514 402618 124546 402854
rect 124782 402618 124866 402854
rect 125102 402618 125134 402854
rect 124514 367174 125134 402618
rect 124514 366938 124546 367174
rect 124782 366938 124866 367174
rect 125102 366938 125134 367174
rect 124514 366854 125134 366938
rect 124514 366618 124546 366854
rect 124782 366618 124866 366854
rect 125102 366618 125134 366854
rect 124514 331174 125134 366618
rect 124514 330938 124546 331174
rect 124782 330938 124866 331174
rect 125102 330938 125134 331174
rect 124514 330854 125134 330938
rect 124514 330618 124546 330854
rect 124782 330618 124866 330854
rect 125102 330618 125134 330854
rect 124514 295174 125134 330618
rect 124514 294938 124546 295174
rect 124782 294938 124866 295174
rect 125102 294938 125134 295174
rect 124514 294854 125134 294938
rect 124514 294618 124546 294854
rect 124782 294618 124866 294854
rect 125102 294618 125134 294854
rect 124514 259174 125134 294618
rect 124514 258938 124546 259174
rect 124782 258938 124866 259174
rect 125102 258938 125134 259174
rect 124514 258854 125134 258938
rect 124514 258618 124546 258854
rect 124782 258618 124866 258854
rect 125102 258618 125134 258854
rect 124514 223174 125134 258618
rect 124514 222938 124546 223174
rect 124782 222938 124866 223174
rect 125102 222938 125134 223174
rect 124514 222854 125134 222938
rect 124514 222618 124546 222854
rect 124782 222618 124866 222854
rect 125102 222618 125134 222854
rect 124514 187174 125134 222618
rect 124514 186938 124546 187174
rect 124782 186938 124866 187174
rect 125102 186938 125134 187174
rect 124514 186854 125134 186938
rect 124514 186618 124546 186854
rect 124782 186618 124866 186854
rect 125102 186618 125134 186854
rect 124514 151174 125134 186618
rect 124514 150938 124546 151174
rect 124782 150938 124866 151174
rect 125102 150938 125134 151174
rect 124514 150854 125134 150938
rect 124514 150618 124546 150854
rect 124782 150618 124866 150854
rect 125102 150618 125134 150854
rect 124514 115174 125134 150618
rect 124514 114938 124546 115174
rect 124782 114938 124866 115174
rect 125102 114938 125134 115174
rect 124514 114854 125134 114938
rect 124514 114618 124546 114854
rect 124782 114618 124866 114854
rect 125102 114618 125134 114854
rect 124514 79174 125134 114618
rect 124514 78938 124546 79174
rect 124782 78938 124866 79174
rect 125102 78938 125134 79174
rect 124514 78854 125134 78938
rect 124514 78618 124546 78854
rect 124782 78618 124866 78854
rect 125102 78618 125134 78854
rect 124514 43174 125134 78618
rect 124514 42938 124546 43174
rect 124782 42938 124866 43174
rect 125102 42938 125134 43174
rect 124514 42854 125134 42938
rect 124514 42618 124546 42854
rect 124782 42618 124866 42854
rect 125102 42618 125134 42854
rect 124514 7174 125134 42618
rect 124514 6938 124546 7174
rect 124782 6938 124866 7174
rect 125102 6938 125134 7174
rect 124514 6854 125134 6938
rect 124514 6618 124546 6854
rect 124782 6618 124866 6854
rect 125102 6618 125134 6854
rect 124514 -2266 125134 6618
rect 124514 -2502 124546 -2266
rect 124782 -2502 124866 -2266
rect 125102 -2502 125134 -2266
rect 124514 -2586 125134 -2502
rect 124514 -2822 124546 -2586
rect 124782 -2822 124866 -2586
rect 125102 -2822 125134 -2586
rect 124514 -3814 125134 -2822
rect 128234 694894 128854 708122
rect 128234 694658 128266 694894
rect 128502 694658 128586 694894
rect 128822 694658 128854 694894
rect 128234 694574 128854 694658
rect 128234 694338 128266 694574
rect 128502 694338 128586 694574
rect 128822 694338 128854 694574
rect 128234 658894 128854 694338
rect 128234 658658 128266 658894
rect 128502 658658 128586 658894
rect 128822 658658 128854 658894
rect 128234 658574 128854 658658
rect 128234 658338 128266 658574
rect 128502 658338 128586 658574
rect 128822 658338 128854 658574
rect 128234 622894 128854 658338
rect 128234 622658 128266 622894
rect 128502 622658 128586 622894
rect 128822 622658 128854 622894
rect 128234 622574 128854 622658
rect 128234 622338 128266 622574
rect 128502 622338 128586 622574
rect 128822 622338 128854 622574
rect 128234 586894 128854 622338
rect 128234 586658 128266 586894
rect 128502 586658 128586 586894
rect 128822 586658 128854 586894
rect 128234 586574 128854 586658
rect 128234 586338 128266 586574
rect 128502 586338 128586 586574
rect 128822 586338 128854 586574
rect 128234 550894 128854 586338
rect 128234 550658 128266 550894
rect 128502 550658 128586 550894
rect 128822 550658 128854 550894
rect 128234 550574 128854 550658
rect 128234 550338 128266 550574
rect 128502 550338 128586 550574
rect 128822 550338 128854 550574
rect 128234 514894 128854 550338
rect 128234 514658 128266 514894
rect 128502 514658 128586 514894
rect 128822 514658 128854 514894
rect 128234 514574 128854 514658
rect 128234 514338 128266 514574
rect 128502 514338 128586 514574
rect 128822 514338 128854 514574
rect 128234 478894 128854 514338
rect 128234 478658 128266 478894
rect 128502 478658 128586 478894
rect 128822 478658 128854 478894
rect 128234 478574 128854 478658
rect 128234 478338 128266 478574
rect 128502 478338 128586 478574
rect 128822 478338 128854 478574
rect 128234 442894 128854 478338
rect 128234 442658 128266 442894
rect 128502 442658 128586 442894
rect 128822 442658 128854 442894
rect 128234 442574 128854 442658
rect 128234 442338 128266 442574
rect 128502 442338 128586 442574
rect 128822 442338 128854 442574
rect 128234 406894 128854 442338
rect 128234 406658 128266 406894
rect 128502 406658 128586 406894
rect 128822 406658 128854 406894
rect 128234 406574 128854 406658
rect 128234 406338 128266 406574
rect 128502 406338 128586 406574
rect 128822 406338 128854 406574
rect 128234 370894 128854 406338
rect 128234 370658 128266 370894
rect 128502 370658 128586 370894
rect 128822 370658 128854 370894
rect 128234 370574 128854 370658
rect 128234 370338 128266 370574
rect 128502 370338 128586 370574
rect 128822 370338 128854 370574
rect 128234 334894 128854 370338
rect 128234 334658 128266 334894
rect 128502 334658 128586 334894
rect 128822 334658 128854 334894
rect 128234 334574 128854 334658
rect 128234 334338 128266 334574
rect 128502 334338 128586 334574
rect 128822 334338 128854 334574
rect 128234 298894 128854 334338
rect 128234 298658 128266 298894
rect 128502 298658 128586 298894
rect 128822 298658 128854 298894
rect 128234 298574 128854 298658
rect 128234 298338 128266 298574
rect 128502 298338 128586 298574
rect 128822 298338 128854 298574
rect 128234 262894 128854 298338
rect 128234 262658 128266 262894
rect 128502 262658 128586 262894
rect 128822 262658 128854 262894
rect 128234 262574 128854 262658
rect 128234 262338 128266 262574
rect 128502 262338 128586 262574
rect 128822 262338 128854 262574
rect 128234 226894 128854 262338
rect 128234 226658 128266 226894
rect 128502 226658 128586 226894
rect 128822 226658 128854 226894
rect 128234 226574 128854 226658
rect 128234 226338 128266 226574
rect 128502 226338 128586 226574
rect 128822 226338 128854 226574
rect 128234 190894 128854 226338
rect 128234 190658 128266 190894
rect 128502 190658 128586 190894
rect 128822 190658 128854 190894
rect 128234 190574 128854 190658
rect 128234 190338 128266 190574
rect 128502 190338 128586 190574
rect 128822 190338 128854 190574
rect 128234 154894 128854 190338
rect 128234 154658 128266 154894
rect 128502 154658 128586 154894
rect 128822 154658 128854 154894
rect 128234 154574 128854 154658
rect 128234 154338 128266 154574
rect 128502 154338 128586 154574
rect 128822 154338 128854 154574
rect 128234 118894 128854 154338
rect 128234 118658 128266 118894
rect 128502 118658 128586 118894
rect 128822 118658 128854 118894
rect 128234 118574 128854 118658
rect 128234 118338 128266 118574
rect 128502 118338 128586 118574
rect 128822 118338 128854 118574
rect 128234 82894 128854 118338
rect 128234 82658 128266 82894
rect 128502 82658 128586 82894
rect 128822 82658 128854 82894
rect 128234 82574 128854 82658
rect 128234 82338 128266 82574
rect 128502 82338 128586 82574
rect 128822 82338 128854 82574
rect 128234 46894 128854 82338
rect 128234 46658 128266 46894
rect 128502 46658 128586 46894
rect 128822 46658 128854 46894
rect 128234 46574 128854 46658
rect 128234 46338 128266 46574
rect 128502 46338 128586 46574
rect 128822 46338 128854 46574
rect 128234 10894 128854 46338
rect 128234 10658 128266 10894
rect 128502 10658 128586 10894
rect 128822 10658 128854 10894
rect 128234 10574 128854 10658
rect 128234 10338 128266 10574
rect 128502 10338 128586 10574
rect 128822 10338 128854 10574
rect 128234 -4186 128854 10338
rect 130794 705798 131414 705830
rect 130794 705562 130826 705798
rect 131062 705562 131146 705798
rect 131382 705562 131414 705798
rect 130794 705478 131414 705562
rect 130794 705242 130826 705478
rect 131062 705242 131146 705478
rect 131382 705242 131414 705478
rect 130794 669454 131414 705242
rect 130794 669218 130826 669454
rect 131062 669218 131146 669454
rect 131382 669218 131414 669454
rect 130794 669134 131414 669218
rect 130794 668898 130826 669134
rect 131062 668898 131146 669134
rect 131382 668898 131414 669134
rect 130794 633454 131414 668898
rect 130794 633218 130826 633454
rect 131062 633218 131146 633454
rect 131382 633218 131414 633454
rect 130794 633134 131414 633218
rect 130794 632898 130826 633134
rect 131062 632898 131146 633134
rect 131382 632898 131414 633134
rect 130794 597454 131414 632898
rect 130794 597218 130826 597454
rect 131062 597218 131146 597454
rect 131382 597218 131414 597454
rect 130794 597134 131414 597218
rect 130794 596898 130826 597134
rect 131062 596898 131146 597134
rect 131382 596898 131414 597134
rect 130794 561454 131414 596898
rect 130794 561218 130826 561454
rect 131062 561218 131146 561454
rect 131382 561218 131414 561454
rect 130794 561134 131414 561218
rect 130794 560898 130826 561134
rect 131062 560898 131146 561134
rect 131382 560898 131414 561134
rect 130794 525454 131414 560898
rect 130794 525218 130826 525454
rect 131062 525218 131146 525454
rect 131382 525218 131414 525454
rect 130794 525134 131414 525218
rect 130794 524898 130826 525134
rect 131062 524898 131146 525134
rect 131382 524898 131414 525134
rect 130794 489454 131414 524898
rect 130794 489218 130826 489454
rect 131062 489218 131146 489454
rect 131382 489218 131414 489454
rect 130794 489134 131414 489218
rect 130794 488898 130826 489134
rect 131062 488898 131146 489134
rect 131382 488898 131414 489134
rect 130794 453454 131414 488898
rect 130794 453218 130826 453454
rect 131062 453218 131146 453454
rect 131382 453218 131414 453454
rect 130794 453134 131414 453218
rect 130794 452898 130826 453134
rect 131062 452898 131146 453134
rect 131382 452898 131414 453134
rect 130794 417454 131414 452898
rect 130794 417218 130826 417454
rect 131062 417218 131146 417454
rect 131382 417218 131414 417454
rect 130794 417134 131414 417218
rect 130794 416898 130826 417134
rect 131062 416898 131146 417134
rect 131382 416898 131414 417134
rect 130794 381454 131414 416898
rect 130794 381218 130826 381454
rect 131062 381218 131146 381454
rect 131382 381218 131414 381454
rect 130794 381134 131414 381218
rect 130794 380898 130826 381134
rect 131062 380898 131146 381134
rect 131382 380898 131414 381134
rect 130794 345454 131414 380898
rect 130794 345218 130826 345454
rect 131062 345218 131146 345454
rect 131382 345218 131414 345454
rect 130794 345134 131414 345218
rect 130794 344898 130826 345134
rect 131062 344898 131146 345134
rect 131382 344898 131414 345134
rect 130794 309454 131414 344898
rect 130794 309218 130826 309454
rect 131062 309218 131146 309454
rect 131382 309218 131414 309454
rect 130794 309134 131414 309218
rect 130794 308898 130826 309134
rect 131062 308898 131146 309134
rect 131382 308898 131414 309134
rect 130794 273454 131414 308898
rect 130794 273218 130826 273454
rect 131062 273218 131146 273454
rect 131382 273218 131414 273454
rect 130794 273134 131414 273218
rect 130794 272898 130826 273134
rect 131062 272898 131146 273134
rect 131382 272898 131414 273134
rect 130794 237454 131414 272898
rect 130794 237218 130826 237454
rect 131062 237218 131146 237454
rect 131382 237218 131414 237454
rect 130794 237134 131414 237218
rect 130794 236898 130826 237134
rect 131062 236898 131146 237134
rect 131382 236898 131414 237134
rect 130794 201454 131414 236898
rect 130794 201218 130826 201454
rect 131062 201218 131146 201454
rect 131382 201218 131414 201454
rect 130794 201134 131414 201218
rect 130794 200898 130826 201134
rect 131062 200898 131146 201134
rect 131382 200898 131414 201134
rect 130794 165454 131414 200898
rect 130794 165218 130826 165454
rect 131062 165218 131146 165454
rect 131382 165218 131414 165454
rect 130794 165134 131414 165218
rect 130794 164898 130826 165134
rect 131062 164898 131146 165134
rect 131382 164898 131414 165134
rect 130794 129454 131414 164898
rect 130794 129218 130826 129454
rect 131062 129218 131146 129454
rect 131382 129218 131414 129454
rect 130794 129134 131414 129218
rect 130794 128898 130826 129134
rect 131062 128898 131146 129134
rect 131382 128898 131414 129134
rect 130794 93454 131414 128898
rect 130794 93218 130826 93454
rect 131062 93218 131146 93454
rect 131382 93218 131414 93454
rect 130794 93134 131414 93218
rect 130794 92898 130826 93134
rect 131062 92898 131146 93134
rect 131382 92898 131414 93134
rect 130794 57454 131414 92898
rect 130794 57218 130826 57454
rect 131062 57218 131146 57454
rect 131382 57218 131414 57454
rect 130794 57134 131414 57218
rect 130794 56898 130826 57134
rect 131062 56898 131146 57134
rect 131382 56898 131414 57134
rect 130794 21454 131414 56898
rect 130794 21218 130826 21454
rect 131062 21218 131146 21454
rect 131382 21218 131414 21454
rect 130794 21134 131414 21218
rect 130794 20898 130826 21134
rect 131062 20898 131146 21134
rect 131382 20898 131414 21134
rect 130794 -1306 131414 20898
rect 130794 -1542 130826 -1306
rect 131062 -1542 131146 -1306
rect 131382 -1542 131414 -1306
rect 130794 -1626 131414 -1542
rect 130794 -1862 130826 -1626
rect 131062 -1862 131146 -1626
rect 131382 -1862 131414 -1626
rect 130794 -1894 131414 -1862
rect 131954 698614 132574 710042
rect 141954 711558 142574 711590
rect 141954 711322 141986 711558
rect 142222 711322 142306 711558
rect 142542 711322 142574 711558
rect 141954 711238 142574 711322
rect 141954 711002 141986 711238
rect 142222 711002 142306 711238
rect 142542 711002 142574 711238
rect 138234 709638 138854 709670
rect 138234 709402 138266 709638
rect 138502 709402 138586 709638
rect 138822 709402 138854 709638
rect 138234 709318 138854 709402
rect 138234 709082 138266 709318
rect 138502 709082 138586 709318
rect 138822 709082 138854 709318
rect 131954 698378 131986 698614
rect 132222 698378 132306 698614
rect 132542 698378 132574 698614
rect 131954 698294 132574 698378
rect 131954 698058 131986 698294
rect 132222 698058 132306 698294
rect 132542 698058 132574 698294
rect 131954 662614 132574 698058
rect 131954 662378 131986 662614
rect 132222 662378 132306 662614
rect 132542 662378 132574 662614
rect 131954 662294 132574 662378
rect 131954 662058 131986 662294
rect 132222 662058 132306 662294
rect 132542 662058 132574 662294
rect 131954 626614 132574 662058
rect 131954 626378 131986 626614
rect 132222 626378 132306 626614
rect 132542 626378 132574 626614
rect 131954 626294 132574 626378
rect 131954 626058 131986 626294
rect 132222 626058 132306 626294
rect 132542 626058 132574 626294
rect 131954 590614 132574 626058
rect 131954 590378 131986 590614
rect 132222 590378 132306 590614
rect 132542 590378 132574 590614
rect 131954 590294 132574 590378
rect 131954 590058 131986 590294
rect 132222 590058 132306 590294
rect 132542 590058 132574 590294
rect 131954 554614 132574 590058
rect 131954 554378 131986 554614
rect 132222 554378 132306 554614
rect 132542 554378 132574 554614
rect 131954 554294 132574 554378
rect 131954 554058 131986 554294
rect 132222 554058 132306 554294
rect 132542 554058 132574 554294
rect 131954 518614 132574 554058
rect 131954 518378 131986 518614
rect 132222 518378 132306 518614
rect 132542 518378 132574 518614
rect 131954 518294 132574 518378
rect 131954 518058 131986 518294
rect 132222 518058 132306 518294
rect 132542 518058 132574 518294
rect 131954 482614 132574 518058
rect 131954 482378 131986 482614
rect 132222 482378 132306 482614
rect 132542 482378 132574 482614
rect 131954 482294 132574 482378
rect 131954 482058 131986 482294
rect 132222 482058 132306 482294
rect 132542 482058 132574 482294
rect 131954 446614 132574 482058
rect 131954 446378 131986 446614
rect 132222 446378 132306 446614
rect 132542 446378 132574 446614
rect 131954 446294 132574 446378
rect 131954 446058 131986 446294
rect 132222 446058 132306 446294
rect 132542 446058 132574 446294
rect 131954 410614 132574 446058
rect 131954 410378 131986 410614
rect 132222 410378 132306 410614
rect 132542 410378 132574 410614
rect 131954 410294 132574 410378
rect 131954 410058 131986 410294
rect 132222 410058 132306 410294
rect 132542 410058 132574 410294
rect 131954 374614 132574 410058
rect 131954 374378 131986 374614
rect 132222 374378 132306 374614
rect 132542 374378 132574 374614
rect 131954 374294 132574 374378
rect 131954 374058 131986 374294
rect 132222 374058 132306 374294
rect 132542 374058 132574 374294
rect 131954 338614 132574 374058
rect 131954 338378 131986 338614
rect 132222 338378 132306 338614
rect 132542 338378 132574 338614
rect 131954 338294 132574 338378
rect 131954 338058 131986 338294
rect 132222 338058 132306 338294
rect 132542 338058 132574 338294
rect 131954 302614 132574 338058
rect 131954 302378 131986 302614
rect 132222 302378 132306 302614
rect 132542 302378 132574 302614
rect 131954 302294 132574 302378
rect 131954 302058 131986 302294
rect 132222 302058 132306 302294
rect 132542 302058 132574 302294
rect 131954 266614 132574 302058
rect 131954 266378 131986 266614
rect 132222 266378 132306 266614
rect 132542 266378 132574 266614
rect 131954 266294 132574 266378
rect 131954 266058 131986 266294
rect 132222 266058 132306 266294
rect 132542 266058 132574 266294
rect 131954 230614 132574 266058
rect 131954 230378 131986 230614
rect 132222 230378 132306 230614
rect 132542 230378 132574 230614
rect 131954 230294 132574 230378
rect 131954 230058 131986 230294
rect 132222 230058 132306 230294
rect 132542 230058 132574 230294
rect 131954 194614 132574 230058
rect 131954 194378 131986 194614
rect 132222 194378 132306 194614
rect 132542 194378 132574 194614
rect 131954 194294 132574 194378
rect 131954 194058 131986 194294
rect 132222 194058 132306 194294
rect 132542 194058 132574 194294
rect 131954 158614 132574 194058
rect 131954 158378 131986 158614
rect 132222 158378 132306 158614
rect 132542 158378 132574 158614
rect 131954 158294 132574 158378
rect 131954 158058 131986 158294
rect 132222 158058 132306 158294
rect 132542 158058 132574 158294
rect 131954 122614 132574 158058
rect 131954 122378 131986 122614
rect 132222 122378 132306 122614
rect 132542 122378 132574 122614
rect 131954 122294 132574 122378
rect 131954 122058 131986 122294
rect 132222 122058 132306 122294
rect 132542 122058 132574 122294
rect 131954 86614 132574 122058
rect 131954 86378 131986 86614
rect 132222 86378 132306 86614
rect 132542 86378 132574 86614
rect 131954 86294 132574 86378
rect 131954 86058 131986 86294
rect 132222 86058 132306 86294
rect 132542 86058 132574 86294
rect 131954 50614 132574 86058
rect 131954 50378 131986 50614
rect 132222 50378 132306 50614
rect 132542 50378 132574 50614
rect 131954 50294 132574 50378
rect 131954 50058 131986 50294
rect 132222 50058 132306 50294
rect 132542 50058 132574 50294
rect 131954 14614 132574 50058
rect 131954 14378 131986 14614
rect 132222 14378 132306 14614
rect 132542 14378 132574 14614
rect 131954 14294 132574 14378
rect 131954 14058 131986 14294
rect 132222 14058 132306 14294
rect 132542 14058 132574 14294
rect 128234 -4422 128266 -4186
rect 128502 -4422 128586 -4186
rect 128822 -4422 128854 -4186
rect 128234 -4506 128854 -4422
rect 128234 -4742 128266 -4506
rect 128502 -4742 128586 -4506
rect 128822 -4742 128854 -4506
rect 128234 -5734 128854 -4742
rect 121954 -7302 121986 -7066
rect 122222 -7302 122306 -7066
rect 122542 -7302 122574 -7066
rect 121954 -7386 122574 -7302
rect 121954 -7622 121986 -7386
rect 122222 -7622 122306 -7386
rect 122542 -7622 122574 -7386
rect 121954 -7654 122574 -7622
rect 131954 -6106 132574 14058
rect 134514 707718 135134 707750
rect 134514 707482 134546 707718
rect 134782 707482 134866 707718
rect 135102 707482 135134 707718
rect 134514 707398 135134 707482
rect 134514 707162 134546 707398
rect 134782 707162 134866 707398
rect 135102 707162 135134 707398
rect 134514 673174 135134 707162
rect 134514 672938 134546 673174
rect 134782 672938 134866 673174
rect 135102 672938 135134 673174
rect 134514 672854 135134 672938
rect 134514 672618 134546 672854
rect 134782 672618 134866 672854
rect 135102 672618 135134 672854
rect 134514 637174 135134 672618
rect 134514 636938 134546 637174
rect 134782 636938 134866 637174
rect 135102 636938 135134 637174
rect 134514 636854 135134 636938
rect 134514 636618 134546 636854
rect 134782 636618 134866 636854
rect 135102 636618 135134 636854
rect 134514 601174 135134 636618
rect 134514 600938 134546 601174
rect 134782 600938 134866 601174
rect 135102 600938 135134 601174
rect 134514 600854 135134 600938
rect 134514 600618 134546 600854
rect 134782 600618 134866 600854
rect 135102 600618 135134 600854
rect 134514 565174 135134 600618
rect 134514 564938 134546 565174
rect 134782 564938 134866 565174
rect 135102 564938 135134 565174
rect 134514 564854 135134 564938
rect 134514 564618 134546 564854
rect 134782 564618 134866 564854
rect 135102 564618 135134 564854
rect 134514 529174 135134 564618
rect 134514 528938 134546 529174
rect 134782 528938 134866 529174
rect 135102 528938 135134 529174
rect 134514 528854 135134 528938
rect 134514 528618 134546 528854
rect 134782 528618 134866 528854
rect 135102 528618 135134 528854
rect 134514 493174 135134 528618
rect 134514 492938 134546 493174
rect 134782 492938 134866 493174
rect 135102 492938 135134 493174
rect 134514 492854 135134 492938
rect 134514 492618 134546 492854
rect 134782 492618 134866 492854
rect 135102 492618 135134 492854
rect 134514 457174 135134 492618
rect 134514 456938 134546 457174
rect 134782 456938 134866 457174
rect 135102 456938 135134 457174
rect 134514 456854 135134 456938
rect 134514 456618 134546 456854
rect 134782 456618 134866 456854
rect 135102 456618 135134 456854
rect 134514 421174 135134 456618
rect 134514 420938 134546 421174
rect 134782 420938 134866 421174
rect 135102 420938 135134 421174
rect 134514 420854 135134 420938
rect 134514 420618 134546 420854
rect 134782 420618 134866 420854
rect 135102 420618 135134 420854
rect 134514 385174 135134 420618
rect 134514 384938 134546 385174
rect 134782 384938 134866 385174
rect 135102 384938 135134 385174
rect 134514 384854 135134 384938
rect 134514 384618 134546 384854
rect 134782 384618 134866 384854
rect 135102 384618 135134 384854
rect 134514 349174 135134 384618
rect 134514 348938 134546 349174
rect 134782 348938 134866 349174
rect 135102 348938 135134 349174
rect 134514 348854 135134 348938
rect 134514 348618 134546 348854
rect 134782 348618 134866 348854
rect 135102 348618 135134 348854
rect 134514 313174 135134 348618
rect 134514 312938 134546 313174
rect 134782 312938 134866 313174
rect 135102 312938 135134 313174
rect 134514 312854 135134 312938
rect 134514 312618 134546 312854
rect 134782 312618 134866 312854
rect 135102 312618 135134 312854
rect 134514 277174 135134 312618
rect 134514 276938 134546 277174
rect 134782 276938 134866 277174
rect 135102 276938 135134 277174
rect 134514 276854 135134 276938
rect 134514 276618 134546 276854
rect 134782 276618 134866 276854
rect 135102 276618 135134 276854
rect 134514 241174 135134 276618
rect 134514 240938 134546 241174
rect 134782 240938 134866 241174
rect 135102 240938 135134 241174
rect 134514 240854 135134 240938
rect 134514 240618 134546 240854
rect 134782 240618 134866 240854
rect 135102 240618 135134 240854
rect 134514 205174 135134 240618
rect 134514 204938 134546 205174
rect 134782 204938 134866 205174
rect 135102 204938 135134 205174
rect 134514 204854 135134 204938
rect 134514 204618 134546 204854
rect 134782 204618 134866 204854
rect 135102 204618 135134 204854
rect 134514 169174 135134 204618
rect 134514 168938 134546 169174
rect 134782 168938 134866 169174
rect 135102 168938 135134 169174
rect 134514 168854 135134 168938
rect 134514 168618 134546 168854
rect 134782 168618 134866 168854
rect 135102 168618 135134 168854
rect 134514 133174 135134 168618
rect 134514 132938 134546 133174
rect 134782 132938 134866 133174
rect 135102 132938 135134 133174
rect 134514 132854 135134 132938
rect 134514 132618 134546 132854
rect 134782 132618 134866 132854
rect 135102 132618 135134 132854
rect 134514 97174 135134 132618
rect 134514 96938 134546 97174
rect 134782 96938 134866 97174
rect 135102 96938 135134 97174
rect 134514 96854 135134 96938
rect 134514 96618 134546 96854
rect 134782 96618 134866 96854
rect 135102 96618 135134 96854
rect 134514 61174 135134 96618
rect 134514 60938 134546 61174
rect 134782 60938 134866 61174
rect 135102 60938 135134 61174
rect 134514 60854 135134 60938
rect 134514 60618 134546 60854
rect 134782 60618 134866 60854
rect 135102 60618 135134 60854
rect 134514 25174 135134 60618
rect 134514 24938 134546 25174
rect 134782 24938 134866 25174
rect 135102 24938 135134 25174
rect 134514 24854 135134 24938
rect 134514 24618 134546 24854
rect 134782 24618 134866 24854
rect 135102 24618 135134 24854
rect 134514 -3226 135134 24618
rect 134514 -3462 134546 -3226
rect 134782 -3462 134866 -3226
rect 135102 -3462 135134 -3226
rect 134514 -3546 135134 -3462
rect 134514 -3782 134546 -3546
rect 134782 -3782 134866 -3546
rect 135102 -3782 135134 -3546
rect 134514 -3814 135134 -3782
rect 138234 676894 138854 709082
rect 138234 676658 138266 676894
rect 138502 676658 138586 676894
rect 138822 676658 138854 676894
rect 138234 676574 138854 676658
rect 138234 676338 138266 676574
rect 138502 676338 138586 676574
rect 138822 676338 138854 676574
rect 138234 640894 138854 676338
rect 138234 640658 138266 640894
rect 138502 640658 138586 640894
rect 138822 640658 138854 640894
rect 138234 640574 138854 640658
rect 138234 640338 138266 640574
rect 138502 640338 138586 640574
rect 138822 640338 138854 640574
rect 138234 604894 138854 640338
rect 138234 604658 138266 604894
rect 138502 604658 138586 604894
rect 138822 604658 138854 604894
rect 138234 604574 138854 604658
rect 138234 604338 138266 604574
rect 138502 604338 138586 604574
rect 138822 604338 138854 604574
rect 138234 568894 138854 604338
rect 138234 568658 138266 568894
rect 138502 568658 138586 568894
rect 138822 568658 138854 568894
rect 138234 568574 138854 568658
rect 138234 568338 138266 568574
rect 138502 568338 138586 568574
rect 138822 568338 138854 568574
rect 138234 532894 138854 568338
rect 138234 532658 138266 532894
rect 138502 532658 138586 532894
rect 138822 532658 138854 532894
rect 138234 532574 138854 532658
rect 138234 532338 138266 532574
rect 138502 532338 138586 532574
rect 138822 532338 138854 532574
rect 138234 496894 138854 532338
rect 138234 496658 138266 496894
rect 138502 496658 138586 496894
rect 138822 496658 138854 496894
rect 138234 496574 138854 496658
rect 138234 496338 138266 496574
rect 138502 496338 138586 496574
rect 138822 496338 138854 496574
rect 138234 460894 138854 496338
rect 138234 460658 138266 460894
rect 138502 460658 138586 460894
rect 138822 460658 138854 460894
rect 138234 460574 138854 460658
rect 138234 460338 138266 460574
rect 138502 460338 138586 460574
rect 138822 460338 138854 460574
rect 138234 424894 138854 460338
rect 138234 424658 138266 424894
rect 138502 424658 138586 424894
rect 138822 424658 138854 424894
rect 138234 424574 138854 424658
rect 138234 424338 138266 424574
rect 138502 424338 138586 424574
rect 138822 424338 138854 424574
rect 138234 388894 138854 424338
rect 138234 388658 138266 388894
rect 138502 388658 138586 388894
rect 138822 388658 138854 388894
rect 138234 388574 138854 388658
rect 138234 388338 138266 388574
rect 138502 388338 138586 388574
rect 138822 388338 138854 388574
rect 138234 352894 138854 388338
rect 138234 352658 138266 352894
rect 138502 352658 138586 352894
rect 138822 352658 138854 352894
rect 138234 352574 138854 352658
rect 138234 352338 138266 352574
rect 138502 352338 138586 352574
rect 138822 352338 138854 352574
rect 138234 316894 138854 352338
rect 138234 316658 138266 316894
rect 138502 316658 138586 316894
rect 138822 316658 138854 316894
rect 138234 316574 138854 316658
rect 138234 316338 138266 316574
rect 138502 316338 138586 316574
rect 138822 316338 138854 316574
rect 138234 280894 138854 316338
rect 138234 280658 138266 280894
rect 138502 280658 138586 280894
rect 138822 280658 138854 280894
rect 138234 280574 138854 280658
rect 138234 280338 138266 280574
rect 138502 280338 138586 280574
rect 138822 280338 138854 280574
rect 138234 244894 138854 280338
rect 138234 244658 138266 244894
rect 138502 244658 138586 244894
rect 138822 244658 138854 244894
rect 138234 244574 138854 244658
rect 138234 244338 138266 244574
rect 138502 244338 138586 244574
rect 138822 244338 138854 244574
rect 138234 208894 138854 244338
rect 138234 208658 138266 208894
rect 138502 208658 138586 208894
rect 138822 208658 138854 208894
rect 138234 208574 138854 208658
rect 138234 208338 138266 208574
rect 138502 208338 138586 208574
rect 138822 208338 138854 208574
rect 138234 172894 138854 208338
rect 138234 172658 138266 172894
rect 138502 172658 138586 172894
rect 138822 172658 138854 172894
rect 138234 172574 138854 172658
rect 138234 172338 138266 172574
rect 138502 172338 138586 172574
rect 138822 172338 138854 172574
rect 138234 136894 138854 172338
rect 138234 136658 138266 136894
rect 138502 136658 138586 136894
rect 138822 136658 138854 136894
rect 138234 136574 138854 136658
rect 138234 136338 138266 136574
rect 138502 136338 138586 136574
rect 138822 136338 138854 136574
rect 138234 100894 138854 136338
rect 138234 100658 138266 100894
rect 138502 100658 138586 100894
rect 138822 100658 138854 100894
rect 138234 100574 138854 100658
rect 138234 100338 138266 100574
rect 138502 100338 138586 100574
rect 138822 100338 138854 100574
rect 138234 64894 138854 100338
rect 138234 64658 138266 64894
rect 138502 64658 138586 64894
rect 138822 64658 138854 64894
rect 138234 64574 138854 64658
rect 138234 64338 138266 64574
rect 138502 64338 138586 64574
rect 138822 64338 138854 64574
rect 138234 28894 138854 64338
rect 138234 28658 138266 28894
rect 138502 28658 138586 28894
rect 138822 28658 138854 28894
rect 138234 28574 138854 28658
rect 138234 28338 138266 28574
rect 138502 28338 138586 28574
rect 138822 28338 138854 28574
rect 138234 -5146 138854 28338
rect 140794 704838 141414 705830
rect 140794 704602 140826 704838
rect 141062 704602 141146 704838
rect 141382 704602 141414 704838
rect 140794 704518 141414 704602
rect 140794 704282 140826 704518
rect 141062 704282 141146 704518
rect 141382 704282 141414 704518
rect 140794 687454 141414 704282
rect 140794 687218 140826 687454
rect 141062 687218 141146 687454
rect 141382 687218 141414 687454
rect 140794 687134 141414 687218
rect 140794 686898 140826 687134
rect 141062 686898 141146 687134
rect 141382 686898 141414 687134
rect 140794 651454 141414 686898
rect 140794 651218 140826 651454
rect 141062 651218 141146 651454
rect 141382 651218 141414 651454
rect 140794 651134 141414 651218
rect 140794 650898 140826 651134
rect 141062 650898 141146 651134
rect 141382 650898 141414 651134
rect 140794 615454 141414 650898
rect 140794 615218 140826 615454
rect 141062 615218 141146 615454
rect 141382 615218 141414 615454
rect 140794 615134 141414 615218
rect 140794 614898 140826 615134
rect 141062 614898 141146 615134
rect 141382 614898 141414 615134
rect 140794 579454 141414 614898
rect 140794 579218 140826 579454
rect 141062 579218 141146 579454
rect 141382 579218 141414 579454
rect 140794 579134 141414 579218
rect 140794 578898 140826 579134
rect 141062 578898 141146 579134
rect 141382 578898 141414 579134
rect 140794 543454 141414 578898
rect 140794 543218 140826 543454
rect 141062 543218 141146 543454
rect 141382 543218 141414 543454
rect 140794 543134 141414 543218
rect 140794 542898 140826 543134
rect 141062 542898 141146 543134
rect 141382 542898 141414 543134
rect 140794 507454 141414 542898
rect 140794 507218 140826 507454
rect 141062 507218 141146 507454
rect 141382 507218 141414 507454
rect 140794 507134 141414 507218
rect 140794 506898 140826 507134
rect 141062 506898 141146 507134
rect 141382 506898 141414 507134
rect 140794 471454 141414 506898
rect 140794 471218 140826 471454
rect 141062 471218 141146 471454
rect 141382 471218 141414 471454
rect 140794 471134 141414 471218
rect 140794 470898 140826 471134
rect 141062 470898 141146 471134
rect 141382 470898 141414 471134
rect 140794 435454 141414 470898
rect 140794 435218 140826 435454
rect 141062 435218 141146 435454
rect 141382 435218 141414 435454
rect 140794 435134 141414 435218
rect 140794 434898 140826 435134
rect 141062 434898 141146 435134
rect 141382 434898 141414 435134
rect 140794 399454 141414 434898
rect 140794 399218 140826 399454
rect 141062 399218 141146 399454
rect 141382 399218 141414 399454
rect 140794 399134 141414 399218
rect 140794 398898 140826 399134
rect 141062 398898 141146 399134
rect 141382 398898 141414 399134
rect 140794 363454 141414 398898
rect 140794 363218 140826 363454
rect 141062 363218 141146 363454
rect 141382 363218 141414 363454
rect 140794 363134 141414 363218
rect 140794 362898 140826 363134
rect 141062 362898 141146 363134
rect 141382 362898 141414 363134
rect 140794 327454 141414 362898
rect 140794 327218 140826 327454
rect 141062 327218 141146 327454
rect 141382 327218 141414 327454
rect 140794 327134 141414 327218
rect 140794 326898 140826 327134
rect 141062 326898 141146 327134
rect 141382 326898 141414 327134
rect 140794 291454 141414 326898
rect 140794 291218 140826 291454
rect 141062 291218 141146 291454
rect 141382 291218 141414 291454
rect 140794 291134 141414 291218
rect 140794 290898 140826 291134
rect 141062 290898 141146 291134
rect 141382 290898 141414 291134
rect 140794 255454 141414 290898
rect 140794 255218 140826 255454
rect 141062 255218 141146 255454
rect 141382 255218 141414 255454
rect 140794 255134 141414 255218
rect 140794 254898 140826 255134
rect 141062 254898 141146 255134
rect 141382 254898 141414 255134
rect 140794 219454 141414 254898
rect 140794 219218 140826 219454
rect 141062 219218 141146 219454
rect 141382 219218 141414 219454
rect 140794 219134 141414 219218
rect 140794 218898 140826 219134
rect 141062 218898 141146 219134
rect 141382 218898 141414 219134
rect 140794 183454 141414 218898
rect 140794 183218 140826 183454
rect 141062 183218 141146 183454
rect 141382 183218 141414 183454
rect 140794 183134 141414 183218
rect 140794 182898 140826 183134
rect 141062 182898 141146 183134
rect 141382 182898 141414 183134
rect 140794 147454 141414 182898
rect 140794 147218 140826 147454
rect 141062 147218 141146 147454
rect 141382 147218 141414 147454
rect 140794 147134 141414 147218
rect 140794 146898 140826 147134
rect 141062 146898 141146 147134
rect 141382 146898 141414 147134
rect 140794 111454 141414 146898
rect 140794 111218 140826 111454
rect 141062 111218 141146 111454
rect 141382 111218 141414 111454
rect 140794 111134 141414 111218
rect 140794 110898 140826 111134
rect 141062 110898 141146 111134
rect 141382 110898 141414 111134
rect 140794 75454 141414 110898
rect 140794 75218 140826 75454
rect 141062 75218 141146 75454
rect 141382 75218 141414 75454
rect 140794 75134 141414 75218
rect 140794 74898 140826 75134
rect 141062 74898 141146 75134
rect 141382 74898 141414 75134
rect 140794 39454 141414 74898
rect 140794 39218 140826 39454
rect 141062 39218 141146 39454
rect 141382 39218 141414 39454
rect 140794 39134 141414 39218
rect 140794 38898 140826 39134
rect 141062 38898 141146 39134
rect 141382 38898 141414 39134
rect 140794 3454 141414 38898
rect 140794 3218 140826 3454
rect 141062 3218 141146 3454
rect 141382 3218 141414 3454
rect 140794 3134 141414 3218
rect 140794 2898 140826 3134
rect 141062 2898 141146 3134
rect 141382 2898 141414 3134
rect 140794 -346 141414 2898
rect 140794 -582 140826 -346
rect 141062 -582 141146 -346
rect 141382 -582 141414 -346
rect 140794 -666 141414 -582
rect 140794 -902 140826 -666
rect 141062 -902 141146 -666
rect 141382 -902 141414 -666
rect 140794 -1894 141414 -902
rect 141954 680614 142574 711002
rect 151954 710598 152574 711590
rect 151954 710362 151986 710598
rect 152222 710362 152306 710598
rect 152542 710362 152574 710598
rect 151954 710278 152574 710362
rect 151954 710042 151986 710278
rect 152222 710042 152306 710278
rect 152542 710042 152574 710278
rect 148234 708678 148854 709670
rect 148234 708442 148266 708678
rect 148502 708442 148586 708678
rect 148822 708442 148854 708678
rect 148234 708358 148854 708442
rect 148234 708122 148266 708358
rect 148502 708122 148586 708358
rect 148822 708122 148854 708358
rect 141954 680378 141986 680614
rect 142222 680378 142306 680614
rect 142542 680378 142574 680614
rect 141954 680294 142574 680378
rect 141954 680058 141986 680294
rect 142222 680058 142306 680294
rect 142542 680058 142574 680294
rect 141954 644614 142574 680058
rect 141954 644378 141986 644614
rect 142222 644378 142306 644614
rect 142542 644378 142574 644614
rect 141954 644294 142574 644378
rect 141954 644058 141986 644294
rect 142222 644058 142306 644294
rect 142542 644058 142574 644294
rect 141954 608614 142574 644058
rect 141954 608378 141986 608614
rect 142222 608378 142306 608614
rect 142542 608378 142574 608614
rect 141954 608294 142574 608378
rect 141954 608058 141986 608294
rect 142222 608058 142306 608294
rect 142542 608058 142574 608294
rect 141954 572614 142574 608058
rect 141954 572378 141986 572614
rect 142222 572378 142306 572614
rect 142542 572378 142574 572614
rect 141954 572294 142574 572378
rect 141954 572058 141986 572294
rect 142222 572058 142306 572294
rect 142542 572058 142574 572294
rect 141954 536614 142574 572058
rect 141954 536378 141986 536614
rect 142222 536378 142306 536614
rect 142542 536378 142574 536614
rect 141954 536294 142574 536378
rect 141954 536058 141986 536294
rect 142222 536058 142306 536294
rect 142542 536058 142574 536294
rect 141954 500614 142574 536058
rect 141954 500378 141986 500614
rect 142222 500378 142306 500614
rect 142542 500378 142574 500614
rect 141954 500294 142574 500378
rect 141954 500058 141986 500294
rect 142222 500058 142306 500294
rect 142542 500058 142574 500294
rect 141954 464614 142574 500058
rect 141954 464378 141986 464614
rect 142222 464378 142306 464614
rect 142542 464378 142574 464614
rect 141954 464294 142574 464378
rect 141954 464058 141986 464294
rect 142222 464058 142306 464294
rect 142542 464058 142574 464294
rect 141954 428614 142574 464058
rect 141954 428378 141986 428614
rect 142222 428378 142306 428614
rect 142542 428378 142574 428614
rect 141954 428294 142574 428378
rect 141954 428058 141986 428294
rect 142222 428058 142306 428294
rect 142542 428058 142574 428294
rect 141954 392614 142574 428058
rect 141954 392378 141986 392614
rect 142222 392378 142306 392614
rect 142542 392378 142574 392614
rect 141954 392294 142574 392378
rect 141954 392058 141986 392294
rect 142222 392058 142306 392294
rect 142542 392058 142574 392294
rect 141954 356614 142574 392058
rect 141954 356378 141986 356614
rect 142222 356378 142306 356614
rect 142542 356378 142574 356614
rect 141954 356294 142574 356378
rect 141954 356058 141986 356294
rect 142222 356058 142306 356294
rect 142542 356058 142574 356294
rect 141954 320614 142574 356058
rect 141954 320378 141986 320614
rect 142222 320378 142306 320614
rect 142542 320378 142574 320614
rect 141954 320294 142574 320378
rect 141954 320058 141986 320294
rect 142222 320058 142306 320294
rect 142542 320058 142574 320294
rect 141954 284614 142574 320058
rect 141954 284378 141986 284614
rect 142222 284378 142306 284614
rect 142542 284378 142574 284614
rect 141954 284294 142574 284378
rect 141954 284058 141986 284294
rect 142222 284058 142306 284294
rect 142542 284058 142574 284294
rect 141954 248614 142574 284058
rect 141954 248378 141986 248614
rect 142222 248378 142306 248614
rect 142542 248378 142574 248614
rect 141954 248294 142574 248378
rect 141954 248058 141986 248294
rect 142222 248058 142306 248294
rect 142542 248058 142574 248294
rect 141954 212614 142574 248058
rect 141954 212378 141986 212614
rect 142222 212378 142306 212614
rect 142542 212378 142574 212614
rect 141954 212294 142574 212378
rect 141954 212058 141986 212294
rect 142222 212058 142306 212294
rect 142542 212058 142574 212294
rect 141954 176614 142574 212058
rect 141954 176378 141986 176614
rect 142222 176378 142306 176614
rect 142542 176378 142574 176614
rect 141954 176294 142574 176378
rect 141954 176058 141986 176294
rect 142222 176058 142306 176294
rect 142542 176058 142574 176294
rect 141954 140614 142574 176058
rect 141954 140378 141986 140614
rect 142222 140378 142306 140614
rect 142542 140378 142574 140614
rect 141954 140294 142574 140378
rect 141954 140058 141986 140294
rect 142222 140058 142306 140294
rect 142542 140058 142574 140294
rect 141954 104614 142574 140058
rect 141954 104378 141986 104614
rect 142222 104378 142306 104614
rect 142542 104378 142574 104614
rect 141954 104294 142574 104378
rect 141954 104058 141986 104294
rect 142222 104058 142306 104294
rect 142542 104058 142574 104294
rect 141954 68614 142574 104058
rect 141954 68378 141986 68614
rect 142222 68378 142306 68614
rect 142542 68378 142574 68614
rect 141954 68294 142574 68378
rect 141954 68058 141986 68294
rect 142222 68058 142306 68294
rect 142542 68058 142574 68294
rect 141954 32614 142574 68058
rect 141954 32378 141986 32614
rect 142222 32378 142306 32614
rect 142542 32378 142574 32614
rect 141954 32294 142574 32378
rect 141954 32058 141986 32294
rect 142222 32058 142306 32294
rect 142542 32058 142574 32294
rect 138234 -5382 138266 -5146
rect 138502 -5382 138586 -5146
rect 138822 -5382 138854 -5146
rect 138234 -5466 138854 -5382
rect 138234 -5702 138266 -5466
rect 138502 -5702 138586 -5466
rect 138822 -5702 138854 -5466
rect 138234 -5734 138854 -5702
rect 131954 -6342 131986 -6106
rect 132222 -6342 132306 -6106
rect 132542 -6342 132574 -6106
rect 131954 -6426 132574 -6342
rect 131954 -6662 131986 -6426
rect 132222 -6662 132306 -6426
rect 132542 -6662 132574 -6426
rect 131954 -7654 132574 -6662
rect 141954 -7066 142574 32058
rect 144514 706758 145134 707750
rect 144514 706522 144546 706758
rect 144782 706522 144866 706758
rect 145102 706522 145134 706758
rect 144514 706438 145134 706522
rect 144514 706202 144546 706438
rect 144782 706202 144866 706438
rect 145102 706202 145134 706438
rect 144514 691174 145134 706202
rect 144514 690938 144546 691174
rect 144782 690938 144866 691174
rect 145102 690938 145134 691174
rect 144514 690854 145134 690938
rect 144514 690618 144546 690854
rect 144782 690618 144866 690854
rect 145102 690618 145134 690854
rect 144514 655174 145134 690618
rect 144514 654938 144546 655174
rect 144782 654938 144866 655174
rect 145102 654938 145134 655174
rect 144514 654854 145134 654938
rect 144514 654618 144546 654854
rect 144782 654618 144866 654854
rect 145102 654618 145134 654854
rect 144514 619174 145134 654618
rect 144514 618938 144546 619174
rect 144782 618938 144866 619174
rect 145102 618938 145134 619174
rect 144514 618854 145134 618938
rect 144514 618618 144546 618854
rect 144782 618618 144866 618854
rect 145102 618618 145134 618854
rect 144514 583174 145134 618618
rect 144514 582938 144546 583174
rect 144782 582938 144866 583174
rect 145102 582938 145134 583174
rect 144514 582854 145134 582938
rect 144514 582618 144546 582854
rect 144782 582618 144866 582854
rect 145102 582618 145134 582854
rect 144514 547174 145134 582618
rect 144514 546938 144546 547174
rect 144782 546938 144866 547174
rect 145102 546938 145134 547174
rect 144514 546854 145134 546938
rect 144514 546618 144546 546854
rect 144782 546618 144866 546854
rect 145102 546618 145134 546854
rect 144514 511174 145134 546618
rect 144514 510938 144546 511174
rect 144782 510938 144866 511174
rect 145102 510938 145134 511174
rect 144514 510854 145134 510938
rect 144514 510618 144546 510854
rect 144782 510618 144866 510854
rect 145102 510618 145134 510854
rect 144514 475174 145134 510618
rect 144514 474938 144546 475174
rect 144782 474938 144866 475174
rect 145102 474938 145134 475174
rect 144514 474854 145134 474938
rect 144514 474618 144546 474854
rect 144782 474618 144866 474854
rect 145102 474618 145134 474854
rect 144514 439174 145134 474618
rect 144514 438938 144546 439174
rect 144782 438938 144866 439174
rect 145102 438938 145134 439174
rect 144514 438854 145134 438938
rect 144514 438618 144546 438854
rect 144782 438618 144866 438854
rect 145102 438618 145134 438854
rect 144514 403174 145134 438618
rect 144514 402938 144546 403174
rect 144782 402938 144866 403174
rect 145102 402938 145134 403174
rect 144514 402854 145134 402938
rect 144514 402618 144546 402854
rect 144782 402618 144866 402854
rect 145102 402618 145134 402854
rect 144514 367174 145134 402618
rect 144514 366938 144546 367174
rect 144782 366938 144866 367174
rect 145102 366938 145134 367174
rect 144514 366854 145134 366938
rect 144514 366618 144546 366854
rect 144782 366618 144866 366854
rect 145102 366618 145134 366854
rect 144514 331174 145134 366618
rect 144514 330938 144546 331174
rect 144782 330938 144866 331174
rect 145102 330938 145134 331174
rect 144514 330854 145134 330938
rect 144514 330618 144546 330854
rect 144782 330618 144866 330854
rect 145102 330618 145134 330854
rect 144514 295174 145134 330618
rect 144514 294938 144546 295174
rect 144782 294938 144866 295174
rect 145102 294938 145134 295174
rect 144514 294854 145134 294938
rect 144514 294618 144546 294854
rect 144782 294618 144866 294854
rect 145102 294618 145134 294854
rect 144514 259174 145134 294618
rect 144514 258938 144546 259174
rect 144782 258938 144866 259174
rect 145102 258938 145134 259174
rect 144514 258854 145134 258938
rect 144514 258618 144546 258854
rect 144782 258618 144866 258854
rect 145102 258618 145134 258854
rect 144514 223174 145134 258618
rect 144514 222938 144546 223174
rect 144782 222938 144866 223174
rect 145102 222938 145134 223174
rect 144514 222854 145134 222938
rect 144514 222618 144546 222854
rect 144782 222618 144866 222854
rect 145102 222618 145134 222854
rect 144514 187174 145134 222618
rect 144514 186938 144546 187174
rect 144782 186938 144866 187174
rect 145102 186938 145134 187174
rect 144514 186854 145134 186938
rect 144514 186618 144546 186854
rect 144782 186618 144866 186854
rect 145102 186618 145134 186854
rect 144514 151174 145134 186618
rect 144514 150938 144546 151174
rect 144782 150938 144866 151174
rect 145102 150938 145134 151174
rect 144514 150854 145134 150938
rect 144514 150618 144546 150854
rect 144782 150618 144866 150854
rect 145102 150618 145134 150854
rect 144514 115174 145134 150618
rect 144514 114938 144546 115174
rect 144782 114938 144866 115174
rect 145102 114938 145134 115174
rect 144514 114854 145134 114938
rect 144514 114618 144546 114854
rect 144782 114618 144866 114854
rect 145102 114618 145134 114854
rect 144514 79174 145134 114618
rect 144514 78938 144546 79174
rect 144782 78938 144866 79174
rect 145102 78938 145134 79174
rect 144514 78854 145134 78938
rect 144514 78618 144546 78854
rect 144782 78618 144866 78854
rect 145102 78618 145134 78854
rect 144514 43174 145134 78618
rect 144514 42938 144546 43174
rect 144782 42938 144866 43174
rect 145102 42938 145134 43174
rect 144514 42854 145134 42938
rect 144514 42618 144546 42854
rect 144782 42618 144866 42854
rect 145102 42618 145134 42854
rect 144514 7174 145134 42618
rect 144514 6938 144546 7174
rect 144782 6938 144866 7174
rect 145102 6938 145134 7174
rect 144514 6854 145134 6938
rect 144514 6618 144546 6854
rect 144782 6618 144866 6854
rect 145102 6618 145134 6854
rect 144514 -2266 145134 6618
rect 144514 -2502 144546 -2266
rect 144782 -2502 144866 -2266
rect 145102 -2502 145134 -2266
rect 144514 -2586 145134 -2502
rect 144514 -2822 144546 -2586
rect 144782 -2822 144866 -2586
rect 145102 -2822 145134 -2586
rect 144514 -3814 145134 -2822
rect 148234 694894 148854 708122
rect 148234 694658 148266 694894
rect 148502 694658 148586 694894
rect 148822 694658 148854 694894
rect 148234 694574 148854 694658
rect 148234 694338 148266 694574
rect 148502 694338 148586 694574
rect 148822 694338 148854 694574
rect 148234 658894 148854 694338
rect 148234 658658 148266 658894
rect 148502 658658 148586 658894
rect 148822 658658 148854 658894
rect 148234 658574 148854 658658
rect 148234 658338 148266 658574
rect 148502 658338 148586 658574
rect 148822 658338 148854 658574
rect 148234 622894 148854 658338
rect 148234 622658 148266 622894
rect 148502 622658 148586 622894
rect 148822 622658 148854 622894
rect 148234 622574 148854 622658
rect 148234 622338 148266 622574
rect 148502 622338 148586 622574
rect 148822 622338 148854 622574
rect 148234 586894 148854 622338
rect 148234 586658 148266 586894
rect 148502 586658 148586 586894
rect 148822 586658 148854 586894
rect 148234 586574 148854 586658
rect 148234 586338 148266 586574
rect 148502 586338 148586 586574
rect 148822 586338 148854 586574
rect 148234 550894 148854 586338
rect 148234 550658 148266 550894
rect 148502 550658 148586 550894
rect 148822 550658 148854 550894
rect 148234 550574 148854 550658
rect 148234 550338 148266 550574
rect 148502 550338 148586 550574
rect 148822 550338 148854 550574
rect 148234 514894 148854 550338
rect 148234 514658 148266 514894
rect 148502 514658 148586 514894
rect 148822 514658 148854 514894
rect 148234 514574 148854 514658
rect 148234 514338 148266 514574
rect 148502 514338 148586 514574
rect 148822 514338 148854 514574
rect 148234 478894 148854 514338
rect 148234 478658 148266 478894
rect 148502 478658 148586 478894
rect 148822 478658 148854 478894
rect 148234 478574 148854 478658
rect 148234 478338 148266 478574
rect 148502 478338 148586 478574
rect 148822 478338 148854 478574
rect 148234 442894 148854 478338
rect 148234 442658 148266 442894
rect 148502 442658 148586 442894
rect 148822 442658 148854 442894
rect 148234 442574 148854 442658
rect 148234 442338 148266 442574
rect 148502 442338 148586 442574
rect 148822 442338 148854 442574
rect 148234 406894 148854 442338
rect 148234 406658 148266 406894
rect 148502 406658 148586 406894
rect 148822 406658 148854 406894
rect 148234 406574 148854 406658
rect 148234 406338 148266 406574
rect 148502 406338 148586 406574
rect 148822 406338 148854 406574
rect 148234 370894 148854 406338
rect 148234 370658 148266 370894
rect 148502 370658 148586 370894
rect 148822 370658 148854 370894
rect 148234 370574 148854 370658
rect 148234 370338 148266 370574
rect 148502 370338 148586 370574
rect 148822 370338 148854 370574
rect 148234 334894 148854 370338
rect 148234 334658 148266 334894
rect 148502 334658 148586 334894
rect 148822 334658 148854 334894
rect 148234 334574 148854 334658
rect 148234 334338 148266 334574
rect 148502 334338 148586 334574
rect 148822 334338 148854 334574
rect 148234 298894 148854 334338
rect 148234 298658 148266 298894
rect 148502 298658 148586 298894
rect 148822 298658 148854 298894
rect 148234 298574 148854 298658
rect 148234 298338 148266 298574
rect 148502 298338 148586 298574
rect 148822 298338 148854 298574
rect 148234 262894 148854 298338
rect 148234 262658 148266 262894
rect 148502 262658 148586 262894
rect 148822 262658 148854 262894
rect 148234 262574 148854 262658
rect 148234 262338 148266 262574
rect 148502 262338 148586 262574
rect 148822 262338 148854 262574
rect 148234 226894 148854 262338
rect 148234 226658 148266 226894
rect 148502 226658 148586 226894
rect 148822 226658 148854 226894
rect 148234 226574 148854 226658
rect 148234 226338 148266 226574
rect 148502 226338 148586 226574
rect 148822 226338 148854 226574
rect 148234 190894 148854 226338
rect 148234 190658 148266 190894
rect 148502 190658 148586 190894
rect 148822 190658 148854 190894
rect 148234 190574 148854 190658
rect 148234 190338 148266 190574
rect 148502 190338 148586 190574
rect 148822 190338 148854 190574
rect 148234 154894 148854 190338
rect 148234 154658 148266 154894
rect 148502 154658 148586 154894
rect 148822 154658 148854 154894
rect 148234 154574 148854 154658
rect 148234 154338 148266 154574
rect 148502 154338 148586 154574
rect 148822 154338 148854 154574
rect 148234 118894 148854 154338
rect 148234 118658 148266 118894
rect 148502 118658 148586 118894
rect 148822 118658 148854 118894
rect 148234 118574 148854 118658
rect 148234 118338 148266 118574
rect 148502 118338 148586 118574
rect 148822 118338 148854 118574
rect 148234 82894 148854 118338
rect 148234 82658 148266 82894
rect 148502 82658 148586 82894
rect 148822 82658 148854 82894
rect 148234 82574 148854 82658
rect 148234 82338 148266 82574
rect 148502 82338 148586 82574
rect 148822 82338 148854 82574
rect 148234 46894 148854 82338
rect 148234 46658 148266 46894
rect 148502 46658 148586 46894
rect 148822 46658 148854 46894
rect 148234 46574 148854 46658
rect 148234 46338 148266 46574
rect 148502 46338 148586 46574
rect 148822 46338 148854 46574
rect 148234 10894 148854 46338
rect 148234 10658 148266 10894
rect 148502 10658 148586 10894
rect 148822 10658 148854 10894
rect 148234 10574 148854 10658
rect 148234 10338 148266 10574
rect 148502 10338 148586 10574
rect 148822 10338 148854 10574
rect 148234 -4186 148854 10338
rect 150794 705798 151414 705830
rect 150794 705562 150826 705798
rect 151062 705562 151146 705798
rect 151382 705562 151414 705798
rect 150794 705478 151414 705562
rect 150794 705242 150826 705478
rect 151062 705242 151146 705478
rect 151382 705242 151414 705478
rect 150794 669454 151414 705242
rect 150794 669218 150826 669454
rect 151062 669218 151146 669454
rect 151382 669218 151414 669454
rect 150794 669134 151414 669218
rect 150794 668898 150826 669134
rect 151062 668898 151146 669134
rect 151382 668898 151414 669134
rect 150794 633454 151414 668898
rect 150794 633218 150826 633454
rect 151062 633218 151146 633454
rect 151382 633218 151414 633454
rect 150794 633134 151414 633218
rect 150794 632898 150826 633134
rect 151062 632898 151146 633134
rect 151382 632898 151414 633134
rect 150794 597454 151414 632898
rect 150794 597218 150826 597454
rect 151062 597218 151146 597454
rect 151382 597218 151414 597454
rect 150794 597134 151414 597218
rect 150794 596898 150826 597134
rect 151062 596898 151146 597134
rect 151382 596898 151414 597134
rect 150794 561454 151414 596898
rect 150794 561218 150826 561454
rect 151062 561218 151146 561454
rect 151382 561218 151414 561454
rect 150794 561134 151414 561218
rect 150794 560898 150826 561134
rect 151062 560898 151146 561134
rect 151382 560898 151414 561134
rect 150794 525454 151414 560898
rect 150794 525218 150826 525454
rect 151062 525218 151146 525454
rect 151382 525218 151414 525454
rect 150794 525134 151414 525218
rect 150794 524898 150826 525134
rect 151062 524898 151146 525134
rect 151382 524898 151414 525134
rect 150794 489454 151414 524898
rect 150794 489218 150826 489454
rect 151062 489218 151146 489454
rect 151382 489218 151414 489454
rect 150794 489134 151414 489218
rect 150794 488898 150826 489134
rect 151062 488898 151146 489134
rect 151382 488898 151414 489134
rect 150794 453454 151414 488898
rect 150794 453218 150826 453454
rect 151062 453218 151146 453454
rect 151382 453218 151414 453454
rect 150794 453134 151414 453218
rect 150794 452898 150826 453134
rect 151062 452898 151146 453134
rect 151382 452898 151414 453134
rect 150794 417454 151414 452898
rect 150794 417218 150826 417454
rect 151062 417218 151146 417454
rect 151382 417218 151414 417454
rect 150794 417134 151414 417218
rect 150794 416898 150826 417134
rect 151062 416898 151146 417134
rect 151382 416898 151414 417134
rect 150794 381454 151414 416898
rect 150794 381218 150826 381454
rect 151062 381218 151146 381454
rect 151382 381218 151414 381454
rect 150794 381134 151414 381218
rect 150794 380898 150826 381134
rect 151062 380898 151146 381134
rect 151382 380898 151414 381134
rect 150794 345454 151414 380898
rect 150794 345218 150826 345454
rect 151062 345218 151146 345454
rect 151382 345218 151414 345454
rect 150794 345134 151414 345218
rect 150794 344898 150826 345134
rect 151062 344898 151146 345134
rect 151382 344898 151414 345134
rect 150794 309454 151414 344898
rect 150794 309218 150826 309454
rect 151062 309218 151146 309454
rect 151382 309218 151414 309454
rect 150794 309134 151414 309218
rect 150794 308898 150826 309134
rect 151062 308898 151146 309134
rect 151382 308898 151414 309134
rect 150794 273454 151414 308898
rect 150794 273218 150826 273454
rect 151062 273218 151146 273454
rect 151382 273218 151414 273454
rect 150794 273134 151414 273218
rect 150794 272898 150826 273134
rect 151062 272898 151146 273134
rect 151382 272898 151414 273134
rect 150794 237454 151414 272898
rect 150794 237218 150826 237454
rect 151062 237218 151146 237454
rect 151382 237218 151414 237454
rect 150794 237134 151414 237218
rect 150794 236898 150826 237134
rect 151062 236898 151146 237134
rect 151382 236898 151414 237134
rect 150794 201454 151414 236898
rect 150794 201218 150826 201454
rect 151062 201218 151146 201454
rect 151382 201218 151414 201454
rect 150794 201134 151414 201218
rect 150794 200898 150826 201134
rect 151062 200898 151146 201134
rect 151382 200898 151414 201134
rect 150794 165454 151414 200898
rect 150794 165218 150826 165454
rect 151062 165218 151146 165454
rect 151382 165218 151414 165454
rect 150794 165134 151414 165218
rect 150794 164898 150826 165134
rect 151062 164898 151146 165134
rect 151382 164898 151414 165134
rect 150794 129454 151414 164898
rect 150794 129218 150826 129454
rect 151062 129218 151146 129454
rect 151382 129218 151414 129454
rect 150794 129134 151414 129218
rect 150794 128898 150826 129134
rect 151062 128898 151146 129134
rect 151382 128898 151414 129134
rect 150794 93454 151414 128898
rect 150794 93218 150826 93454
rect 151062 93218 151146 93454
rect 151382 93218 151414 93454
rect 150794 93134 151414 93218
rect 150794 92898 150826 93134
rect 151062 92898 151146 93134
rect 151382 92898 151414 93134
rect 150794 57454 151414 92898
rect 150794 57218 150826 57454
rect 151062 57218 151146 57454
rect 151382 57218 151414 57454
rect 150794 57134 151414 57218
rect 150794 56898 150826 57134
rect 151062 56898 151146 57134
rect 151382 56898 151414 57134
rect 150794 21454 151414 56898
rect 150794 21218 150826 21454
rect 151062 21218 151146 21454
rect 151382 21218 151414 21454
rect 150794 21134 151414 21218
rect 150794 20898 150826 21134
rect 151062 20898 151146 21134
rect 151382 20898 151414 21134
rect 150794 -1306 151414 20898
rect 150794 -1542 150826 -1306
rect 151062 -1542 151146 -1306
rect 151382 -1542 151414 -1306
rect 150794 -1626 151414 -1542
rect 150794 -1862 150826 -1626
rect 151062 -1862 151146 -1626
rect 151382 -1862 151414 -1626
rect 150794 -1894 151414 -1862
rect 151954 698614 152574 710042
rect 161954 711558 162574 711590
rect 161954 711322 161986 711558
rect 162222 711322 162306 711558
rect 162542 711322 162574 711558
rect 161954 711238 162574 711322
rect 161954 711002 161986 711238
rect 162222 711002 162306 711238
rect 162542 711002 162574 711238
rect 158234 709638 158854 709670
rect 158234 709402 158266 709638
rect 158502 709402 158586 709638
rect 158822 709402 158854 709638
rect 158234 709318 158854 709402
rect 158234 709082 158266 709318
rect 158502 709082 158586 709318
rect 158822 709082 158854 709318
rect 151954 698378 151986 698614
rect 152222 698378 152306 698614
rect 152542 698378 152574 698614
rect 151954 698294 152574 698378
rect 151954 698058 151986 698294
rect 152222 698058 152306 698294
rect 152542 698058 152574 698294
rect 151954 662614 152574 698058
rect 151954 662378 151986 662614
rect 152222 662378 152306 662614
rect 152542 662378 152574 662614
rect 151954 662294 152574 662378
rect 151954 662058 151986 662294
rect 152222 662058 152306 662294
rect 152542 662058 152574 662294
rect 151954 626614 152574 662058
rect 151954 626378 151986 626614
rect 152222 626378 152306 626614
rect 152542 626378 152574 626614
rect 151954 626294 152574 626378
rect 151954 626058 151986 626294
rect 152222 626058 152306 626294
rect 152542 626058 152574 626294
rect 151954 590614 152574 626058
rect 151954 590378 151986 590614
rect 152222 590378 152306 590614
rect 152542 590378 152574 590614
rect 151954 590294 152574 590378
rect 151954 590058 151986 590294
rect 152222 590058 152306 590294
rect 152542 590058 152574 590294
rect 151954 554614 152574 590058
rect 151954 554378 151986 554614
rect 152222 554378 152306 554614
rect 152542 554378 152574 554614
rect 151954 554294 152574 554378
rect 151954 554058 151986 554294
rect 152222 554058 152306 554294
rect 152542 554058 152574 554294
rect 151954 518614 152574 554058
rect 151954 518378 151986 518614
rect 152222 518378 152306 518614
rect 152542 518378 152574 518614
rect 151954 518294 152574 518378
rect 151954 518058 151986 518294
rect 152222 518058 152306 518294
rect 152542 518058 152574 518294
rect 151954 482614 152574 518058
rect 151954 482378 151986 482614
rect 152222 482378 152306 482614
rect 152542 482378 152574 482614
rect 151954 482294 152574 482378
rect 151954 482058 151986 482294
rect 152222 482058 152306 482294
rect 152542 482058 152574 482294
rect 151954 446614 152574 482058
rect 151954 446378 151986 446614
rect 152222 446378 152306 446614
rect 152542 446378 152574 446614
rect 151954 446294 152574 446378
rect 151954 446058 151986 446294
rect 152222 446058 152306 446294
rect 152542 446058 152574 446294
rect 151954 410614 152574 446058
rect 151954 410378 151986 410614
rect 152222 410378 152306 410614
rect 152542 410378 152574 410614
rect 151954 410294 152574 410378
rect 151954 410058 151986 410294
rect 152222 410058 152306 410294
rect 152542 410058 152574 410294
rect 151954 374614 152574 410058
rect 151954 374378 151986 374614
rect 152222 374378 152306 374614
rect 152542 374378 152574 374614
rect 151954 374294 152574 374378
rect 151954 374058 151986 374294
rect 152222 374058 152306 374294
rect 152542 374058 152574 374294
rect 151954 338614 152574 374058
rect 151954 338378 151986 338614
rect 152222 338378 152306 338614
rect 152542 338378 152574 338614
rect 151954 338294 152574 338378
rect 151954 338058 151986 338294
rect 152222 338058 152306 338294
rect 152542 338058 152574 338294
rect 151954 302614 152574 338058
rect 151954 302378 151986 302614
rect 152222 302378 152306 302614
rect 152542 302378 152574 302614
rect 151954 302294 152574 302378
rect 151954 302058 151986 302294
rect 152222 302058 152306 302294
rect 152542 302058 152574 302294
rect 151954 266614 152574 302058
rect 151954 266378 151986 266614
rect 152222 266378 152306 266614
rect 152542 266378 152574 266614
rect 151954 266294 152574 266378
rect 151954 266058 151986 266294
rect 152222 266058 152306 266294
rect 152542 266058 152574 266294
rect 151954 230614 152574 266058
rect 151954 230378 151986 230614
rect 152222 230378 152306 230614
rect 152542 230378 152574 230614
rect 151954 230294 152574 230378
rect 151954 230058 151986 230294
rect 152222 230058 152306 230294
rect 152542 230058 152574 230294
rect 151954 194614 152574 230058
rect 151954 194378 151986 194614
rect 152222 194378 152306 194614
rect 152542 194378 152574 194614
rect 151954 194294 152574 194378
rect 151954 194058 151986 194294
rect 152222 194058 152306 194294
rect 152542 194058 152574 194294
rect 151954 158614 152574 194058
rect 151954 158378 151986 158614
rect 152222 158378 152306 158614
rect 152542 158378 152574 158614
rect 151954 158294 152574 158378
rect 151954 158058 151986 158294
rect 152222 158058 152306 158294
rect 152542 158058 152574 158294
rect 151954 122614 152574 158058
rect 151954 122378 151986 122614
rect 152222 122378 152306 122614
rect 152542 122378 152574 122614
rect 151954 122294 152574 122378
rect 151954 122058 151986 122294
rect 152222 122058 152306 122294
rect 152542 122058 152574 122294
rect 151954 86614 152574 122058
rect 151954 86378 151986 86614
rect 152222 86378 152306 86614
rect 152542 86378 152574 86614
rect 151954 86294 152574 86378
rect 151954 86058 151986 86294
rect 152222 86058 152306 86294
rect 152542 86058 152574 86294
rect 151954 50614 152574 86058
rect 151954 50378 151986 50614
rect 152222 50378 152306 50614
rect 152542 50378 152574 50614
rect 151954 50294 152574 50378
rect 151954 50058 151986 50294
rect 152222 50058 152306 50294
rect 152542 50058 152574 50294
rect 151954 14614 152574 50058
rect 151954 14378 151986 14614
rect 152222 14378 152306 14614
rect 152542 14378 152574 14614
rect 151954 14294 152574 14378
rect 151954 14058 151986 14294
rect 152222 14058 152306 14294
rect 152542 14058 152574 14294
rect 148234 -4422 148266 -4186
rect 148502 -4422 148586 -4186
rect 148822 -4422 148854 -4186
rect 148234 -4506 148854 -4422
rect 148234 -4742 148266 -4506
rect 148502 -4742 148586 -4506
rect 148822 -4742 148854 -4506
rect 148234 -5734 148854 -4742
rect 141954 -7302 141986 -7066
rect 142222 -7302 142306 -7066
rect 142542 -7302 142574 -7066
rect 141954 -7386 142574 -7302
rect 141954 -7622 141986 -7386
rect 142222 -7622 142306 -7386
rect 142542 -7622 142574 -7386
rect 141954 -7654 142574 -7622
rect 151954 -6106 152574 14058
rect 154514 707718 155134 707750
rect 154514 707482 154546 707718
rect 154782 707482 154866 707718
rect 155102 707482 155134 707718
rect 154514 707398 155134 707482
rect 154514 707162 154546 707398
rect 154782 707162 154866 707398
rect 155102 707162 155134 707398
rect 154514 673174 155134 707162
rect 154514 672938 154546 673174
rect 154782 672938 154866 673174
rect 155102 672938 155134 673174
rect 154514 672854 155134 672938
rect 154514 672618 154546 672854
rect 154782 672618 154866 672854
rect 155102 672618 155134 672854
rect 154514 637174 155134 672618
rect 154514 636938 154546 637174
rect 154782 636938 154866 637174
rect 155102 636938 155134 637174
rect 154514 636854 155134 636938
rect 154514 636618 154546 636854
rect 154782 636618 154866 636854
rect 155102 636618 155134 636854
rect 154514 601174 155134 636618
rect 154514 600938 154546 601174
rect 154782 600938 154866 601174
rect 155102 600938 155134 601174
rect 154514 600854 155134 600938
rect 154514 600618 154546 600854
rect 154782 600618 154866 600854
rect 155102 600618 155134 600854
rect 154514 565174 155134 600618
rect 154514 564938 154546 565174
rect 154782 564938 154866 565174
rect 155102 564938 155134 565174
rect 154514 564854 155134 564938
rect 154514 564618 154546 564854
rect 154782 564618 154866 564854
rect 155102 564618 155134 564854
rect 154514 529174 155134 564618
rect 154514 528938 154546 529174
rect 154782 528938 154866 529174
rect 155102 528938 155134 529174
rect 154514 528854 155134 528938
rect 154514 528618 154546 528854
rect 154782 528618 154866 528854
rect 155102 528618 155134 528854
rect 154514 493174 155134 528618
rect 154514 492938 154546 493174
rect 154782 492938 154866 493174
rect 155102 492938 155134 493174
rect 154514 492854 155134 492938
rect 154514 492618 154546 492854
rect 154782 492618 154866 492854
rect 155102 492618 155134 492854
rect 154514 457174 155134 492618
rect 154514 456938 154546 457174
rect 154782 456938 154866 457174
rect 155102 456938 155134 457174
rect 154514 456854 155134 456938
rect 154514 456618 154546 456854
rect 154782 456618 154866 456854
rect 155102 456618 155134 456854
rect 154514 421174 155134 456618
rect 154514 420938 154546 421174
rect 154782 420938 154866 421174
rect 155102 420938 155134 421174
rect 154514 420854 155134 420938
rect 154514 420618 154546 420854
rect 154782 420618 154866 420854
rect 155102 420618 155134 420854
rect 154514 385174 155134 420618
rect 154514 384938 154546 385174
rect 154782 384938 154866 385174
rect 155102 384938 155134 385174
rect 154514 384854 155134 384938
rect 154514 384618 154546 384854
rect 154782 384618 154866 384854
rect 155102 384618 155134 384854
rect 154514 349174 155134 384618
rect 154514 348938 154546 349174
rect 154782 348938 154866 349174
rect 155102 348938 155134 349174
rect 154514 348854 155134 348938
rect 154514 348618 154546 348854
rect 154782 348618 154866 348854
rect 155102 348618 155134 348854
rect 154514 313174 155134 348618
rect 154514 312938 154546 313174
rect 154782 312938 154866 313174
rect 155102 312938 155134 313174
rect 154514 312854 155134 312938
rect 154514 312618 154546 312854
rect 154782 312618 154866 312854
rect 155102 312618 155134 312854
rect 154514 277174 155134 312618
rect 154514 276938 154546 277174
rect 154782 276938 154866 277174
rect 155102 276938 155134 277174
rect 154514 276854 155134 276938
rect 154514 276618 154546 276854
rect 154782 276618 154866 276854
rect 155102 276618 155134 276854
rect 154514 241174 155134 276618
rect 154514 240938 154546 241174
rect 154782 240938 154866 241174
rect 155102 240938 155134 241174
rect 154514 240854 155134 240938
rect 154514 240618 154546 240854
rect 154782 240618 154866 240854
rect 155102 240618 155134 240854
rect 154514 205174 155134 240618
rect 154514 204938 154546 205174
rect 154782 204938 154866 205174
rect 155102 204938 155134 205174
rect 154514 204854 155134 204938
rect 154514 204618 154546 204854
rect 154782 204618 154866 204854
rect 155102 204618 155134 204854
rect 154514 169174 155134 204618
rect 154514 168938 154546 169174
rect 154782 168938 154866 169174
rect 155102 168938 155134 169174
rect 154514 168854 155134 168938
rect 154514 168618 154546 168854
rect 154782 168618 154866 168854
rect 155102 168618 155134 168854
rect 154514 133174 155134 168618
rect 154514 132938 154546 133174
rect 154782 132938 154866 133174
rect 155102 132938 155134 133174
rect 154514 132854 155134 132938
rect 154514 132618 154546 132854
rect 154782 132618 154866 132854
rect 155102 132618 155134 132854
rect 154514 97174 155134 132618
rect 154514 96938 154546 97174
rect 154782 96938 154866 97174
rect 155102 96938 155134 97174
rect 154514 96854 155134 96938
rect 154514 96618 154546 96854
rect 154782 96618 154866 96854
rect 155102 96618 155134 96854
rect 154514 61174 155134 96618
rect 154514 60938 154546 61174
rect 154782 60938 154866 61174
rect 155102 60938 155134 61174
rect 154514 60854 155134 60938
rect 154514 60618 154546 60854
rect 154782 60618 154866 60854
rect 155102 60618 155134 60854
rect 154514 25174 155134 60618
rect 154514 24938 154546 25174
rect 154782 24938 154866 25174
rect 155102 24938 155134 25174
rect 154514 24854 155134 24938
rect 154514 24618 154546 24854
rect 154782 24618 154866 24854
rect 155102 24618 155134 24854
rect 154514 -3226 155134 24618
rect 154514 -3462 154546 -3226
rect 154782 -3462 154866 -3226
rect 155102 -3462 155134 -3226
rect 154514 -3546 155134 -3462
rect 154514 -3782 154546 -3546
rect 154782 -3782 154866 -3546
rect 155102 -3782 155134 -3546
rect 154514 -3814 155134 -3782
rect 158234 676894 158854 709082
rect 158234 676658 158266 676894
rect 158502 676658 158586 676894
rect 158822 676658 158854 676894
rect 158234 676574 158854 676658
rect 158234 676338 158266 676574
rect 158502 676338 158586 676574
rect 158822 676338 158854 676574
rect 158234 640894 158854 676338
rect 158234 640658 158266 640894
rect 158502 640658 158586 640894
rect 158822 640658 158854 640894
rect 158234 640574 158854 640658
rect 158234 640338 158266 640574
rect 158502 640338 158586 640574
rect 158822 640338 158854 640574
rect 158234 604894 158854 640338
rect 158234 604658 158266 604894
rect 158502 604658 158586 604894
rect 158822 604658 158854 604894
rect 158234 604574 158854 604658
rect 158234 604338 158266 604574
rect 158502 604338 158586 604574
rect 158822 604338 158854 604574
rect 158234 568894 158854 604338
rect 158234 568658 158266 568894
rect 158502 568658 158586 568894
rect 158822 568658 158854 568894
rect 158234 568574 158854 568658
rect 158234 568338 158266 568574
rect 158502 568338 158586 568574
rect 158822 568338 158854 568574
rect 158234 532894 158854 568338
rect 158234 532658 158266 532894
rect 158502 532658 158586 532894
rect 158822 532658 158854 532894
rect 158234 532574 158854 532658
rect 158234 532338 158266 532574
rect 158502 532338 158586 532574
rect 158822 532338 158854 532574
rect 158234 496894 158854 532338
rect 158234 496658 158266 496894
rect 158502 496658 158586 496894
rect 158822 496658 158854 496894
rect 158234 496574 158854 496658
rect 158234 496338 158266 496574
rect 158502 496338 158586 496574
rect 158822 496338 158854 496574
rect 158234 460894 158854 496338
rect 158234 460658 158266 460894
rect 158502 460658 158586 460894
rect 158822 460658 158854 460894
rect 158234 460574 158854 460658
rect 158234 460338 158266 460574
rect 158502 460338 158586 460574
rect 158822 460338 158854 460574
rect 158234 424894 158854 460338
rect 158234 424658 158266 424894
rect 158502 424658 158586 424894
rect 158822 424658 158854 424894
rect 158234 424574 158854 424658
rect 158234 424338 158266 424574
rect 158502 424338 158586 424574
rect 158822 424338 158854 424574
rect 158234 388894 158854 424338
rect 158234 388658 158266 388894
rect 158502 388658 158586 388894
rect 158822 388658 158854 388894
rect 158234 388574 158854 388658
rect 158234 388338 158266 388574
rect 158502 388338 158586 388574
rect 158822 388338 158854 388574
rect 158234 352894 158854 388338
rect 158234 352658 158266 352894
rect 158502 352658 158586 352894
rect 158822 352658 158854 352894
rect 158234 352574 158854 352658
rect 158234 352338 158266 352574
rect 158502 352338 158586 352574
rect 158822 352338 158854 352574
rect 158234 316894 158854 352338
rect 158234 316658 158266 316894
rect 158502 316658 158586 316894
rect 158822 316658 158854 316894
rect 158234 316574 158854 316658
rect 158234 316338 158266 316574
rect 158502 316338 158586 316574
rect 158822 316338 158854 316574
rect 158234 280894 158854 316338
rect 158234 280658 158266 280894
rect 158502 280658 158586 280894
rect 158822 280658 158854 280894
rect 158234 280574 158854 280658
rect 158234 280338 158266 280574
rect 158502 280338 158586 280574
rect 158822 280338 158854 280574
rect 158234 244894 158854 280338
rect 158234 244658 158266 244894
rect 158502 244658 158586 244894
rect 158822 244658 158854 244894
rect 158234 244574 158854 244658
rect 158234 244338 158266 244574
rect 158502 244338 158586 244574
rect 158822 244338 158854 244574
rect 158234 208894 158854 244338
rect 158234 208658 158266 208894
rect 158502 208658 158586 208894
rect 158822 208658 158854 208894
rect 158234 208574 158854 208658
rect 158234 208338 158266 208574
rect 158502 208338 158586 208574
rect 158822 208338 158854 208574
rect 158234 172894 158854 208338
rect 158234 172658 158266 172894
rect 158502 172658 158586 172894
rect 158822 172658 158854 172894
rect 158234 172574 158854 172658
rect 158234 172338 158266 172574
rect 158502 172338 158586 172574
rect 158822 172338 158854 172574
rect 158234 136894 158854 172338
rect 158234 136658 158266 136894
rect 158502 136658 158586 136894
rect 158822 136658 158854 136894
rect 158234 136574 158854 136658
rect 158234 136338 158266 136574
rect 158502 136338 158586 136574
rect 158822 136338 158854 136574
rect 158234 100894 158854 136338
rect 158234 100658 158266 100894
rect 158502 100658 158586 100894
rect 158822 100658 158854 100894
rect 158234 100574 158854 100658
rect 158234 100338 158266 100574
rect 158502 100338 158586 100574
rect 158822 100338 158854 100574
rect 158234 64894 158854 100338
rect 158234 64658 158266 64894
rect 158502 64658 158586 64894
rect 158822 64658 158854 64894
rect 158234 64574 158854 64658
rect 158234 64338 158266 64574
rect 158502 64338 158586 64574
rect 158822 64338 158854 64574
rect 158234 28894 158854 64338
rect 158234 28658 158266 28894
rect 158502 28658 158586 28894
rect 158822 28658 158854 28894
rect 158234 28574 158854 28658
rect 158234 28338 158266 28574
rect 158502 28338 158586 28574
rect 158822 28338 158854 28574
rect 158234 -5146 158854 28338
rect 160794 704838 161414 705830
rect 160794 704602 160826 704838
rect 161062 704602 161146 704838
rect 161382 704602 161414 704838
rect 160794 704518 161414 704602
rect 160794 704282 160826 704518
rect 161062 704282 161146 704518
rect 161382 704282 161414 704518
rect 160794 687454 161414 704282
rect 160794 687218 160826 687454
rect 161062 687218 161146 687454
rect 161382 687218 161414 687454
rect 160794 687134 161414 687218
rect 160794 686898 160826 687134
rect 161062 686898 161146 687134
rect 161382 686898 161414 687134
rect 160794 651454 161414 686898
rect 160794 651218 160826 651454
rect 161062 651218 161146 651454
rect 161382 651218 161414 651454
rect 160794 651134 161414 651218
rect 160794 650898 160826 651134
rect 161062 650898 161146 651134
rect 161382 650898 161414 651134
rect 160794 615454 161414 650898
rect 160794 615218 160826 615454
rect 161062 615218 161146 615454
rect 161382 615218 161414 615454
rect 160794 615134 161414 615218
rect 160794 614898 160826 615134
rect 161062 614898 161146 615134
rect 161382 614898 161414 615134
rect 160794 579454 161414 614898
rect 160794 579218 160826 579454
rect 161062 579218 161146 579454
rect 161382 579218 161414 579454
rect 160794 579134 161414 579218
rect 160794 578898 160826 579134
rect 161062 578898 161146 579134
rect 161382 578898 161414 579134
rect 160794 543454 161414 578898
rect 160794 543218 160826 543454
rect 161062 543218 161146 543454
rect 161382 543218 161414 543454
rect 160794 543134 161414 543218
rect 160794 542898 160826 543134
rect 161062 542898 161146 543134
rect 161382 542898 161414 543134
rect 160794 507454 161414 542898
rect 160794 507218 160826 507454
rect 161062 507218 161146 507454
rect 161382 507218 161414 507454
rect 160794 507134 161414 507218
rect 160794 506898 160826 507134
rect 161062 506898 161146 507134
rect 161382 506898 161414 507134
rect 160794 471454 161414 506898
rect 160794 471218 160826 471454
rect 161062 471218 161146 471454
rect 161382 471218 161414 471454
rect 160794 471134 161414 471218
rect 160794 470898 160826 471134
rect 161062 470898 161146 471134
rect 161382 470898 161414 471134
rect 160794 435454 161414 470898
rect 160794 435218 160826 435454
rect 161062 435218 161146 435454
rect 161382 435218 161414 435454
rect 160794 435134 161414 435218
rect 160794 434898 160826 435134
rect 161062 434898 161146 435134
rect 161382 434898 161414 435134
rect 160794 399454 161414 434898
rect 160794 399218 160826 399454
rect 161062 399218 161146 399454
rect 161382 399218 161414 399454
rect 160794 399134 161414 399218
rect 160794 398898 160826 399134
rect 161062 398898 161146 399134
rect 161382 398898 161414 399134
rect 160794 363454 161414 398898
rect 160794 363218 160826 363454
rect 161062 363218 161146 363454
rect 161382 363218 161414 363454
rect 160794 363134 161414 363218
rect 160794 362898 160826 363134
rect 161062 362898 161146 363134
rect 161382 362898 161414 363134
rect 160794 327454 161414 362898
rect 160794 327218 160826 327454
rect 161062 327218 161146 327454
rect 161382 327218 161414 327454
rect 160794 327134 161414 327218
rect 160794 326898 160826 327134
rect 161062 326898 161146 327134
rect 161382 326898 161414 327134
rect 160794 291454 161414 326898
rect 160794 291218 160826 291454
rect 161062 291218 161146 291454
rect 161382 291218 161414 291454
rect 160794 291134 161414 291218
rect 160794 290898 160826 291134
rect 161062 290898 161146 291134
rect 161382 290898 161414 291134
rect 160794 255454 161414 290898
rect 160794 255218 160826 255454
rect 161062 255218 161146 255454
rect 161382 255218 161414 255454
rect 160794 255134 161414 255218
rect 160794 254898 160826 255134
rect 161062 254898 161146 255134
rect 161382 254898 161414 255134
rect 160794 219454 161414 254898
rect 160794 219218 160826 219454
rect 161062 219218 161146 219454
rect 161382 219218 161414 219454
rect 160794 219134 161414 219218
rect 160794 218898 160826 219134
rect 161062 218898 161146 219134
rect 161382 218898 161414 219134
rect 160794 183454 161414 218898
rect 160794 183218 160826 183454
rect 161062 183218 161146 183454
rect 161382 183218 161414 183454
rect 160794 183134 161414 183218
rect 160794 182898 160826 183134
rect 161062 182898 161146 183134
rect 161382 182898 161414 183134
rect 160794 147454 161414 182898
rect 160794 147218 160826 147454
rect 161062 147218 161146 147454
rect 161382 147218 161414 147454
rect 160794 147134 161414 147218
rect 160794 146898 160826 147134
rect 161062 146898 161146 147134
rect 161382 146898 161414 147134
rect 160794 111454 161414 146898
rect 160794 111218 160826 111454
rect 161062 111218 161146 111454
rect 161382 111218 161414 111454
rect 160794 111134 161414 111218
rect 160794 110898 160826 111134
rect 161062 110898 161146 111134
rect 161382 110898 161414 111134
rect 160794 75454 161414 110898
rect 160794 75218 160826 75454
rect 161062 75218 161146 75454
rect 161382 75218 161414 75454
rect 160794 75134 161414 75218
rect 160794 74898 160826 75134
rect 161062 74898 161146 75134
rect 161382 74898 161414 75134
rect 160794 39454 161414 74898
rect 160794 39218 160826 39454
rect 161062 39218 161146 39454
rect 161382 39218 161414 39454
rect 160794 39134 161414 39218
rect 160794 38898 160826 39134
rect 161062 38898 161146 39134
rect 161382 38898 161414 39134
rect 160794 3454 161414 38898
rect 160794 3218 160826 3454
rect 161062 3218 161146 3454
rect 161382 3218 161414 3454
rect 160794 3134 161414 3218
rect 160794 2898 160826 3134
rect 161062 2898 161146 3134
rect 161382 2898 161414 3134
rect 160794 -346 161414 2898
rect 160794 -582 160826 -346
rect 161062 -582 161146 -346
rect 161382 -582 161414 -346
rect 160794 -666 161414 -582
rect 160794 -902 160826 -666
rect 161062 -902 161146 -666
rect 161382 -902 161414 -666
rect 160794 -1894 161414 -902
rect 161954 680614 162574 711002
rect 171954 710598 172574 711590
rect 171954 710362 171986 710598
rect 172222 710362 172306 710598
rect 172542 710362 172574 710598
rect 171954 710278 172574 710362
rect 171954 710042 171986 710278
rect 172222 710042 172306 710278
rect 172542 710042 172574 710278
rect 168234 708678 168854 709670
rect 168234 708442 168266 708678
rect 168502 708442 168586 708678
rect 168822 708442 168854 708678
rect 168234 708358 168854 708442
rect 168234 708122 168266 708358
rect 168502 708122 168586 708358
rect 168822 708122 168854 708358
rect 161954 680378 161986 680614
rect 162222 680378 162306 680614
rect 162542 680378 162574 680614
rect 161954 680294 162574 680378
rect 161954 680058 161986 680294
rect 162222 680058 162306 680294
rect 162542 680058 162574 680294
rect 161954 644614 162574 680058
rect 161954 644378 161986 644614
rect 162222 644378 162306 644614
rect 162542 644378 162574 644614
rect 161954 644294 162574 644378
rect 161954 644058 161986 644294
rect 162222 644058 162306 644294
rect 162542 644058 162574 644294
rect 161954 608614 162574 644058
rect 161954 608378 161986 608614
rect 162222 608378 162306 608614
rect 162542 608378 162574 608614
rect 161954 608294 162574 608378
rect 161954 608058 161986 608294
rect 162222 608058 162306 608294
rect 162542 608058 162574 608294
rect 161954 572614 162574 608058
rect 161954 572378 161986 572614
rect 162222 572378 162306 572614
rect 162542 572378 162574 572614
rect 161954 572294 162574 572378
rect 161954 572058 161986 572294
rect 162222 572058 162306 572294
rect 162542 572058 162574 572294
rect 161954 536614 162574 572058
rect 161954 536378 161986 536614
rect 162222 536378 162306 536614
rect 162542 536378 162574 536614
rect 161954 536294 162574 536378
rect 161954 536058 161986 536294
rect 162222 536058 162306 536294
rect 162542 536058 162574 536294
rect 161954 500614 162574 536058
rect 161954 500378 161986 500614
rect 162222 500378 162306 500614
rect 162542 500378 162574 500614
rect 161954 500294 162574 500378
rect 161954 500058 161986 500294
rect 162222 500058 162306 500294
rect 162542 500058 162574 500294
rect 161954 464614 162574 500058
rect 161954 464378 161986 464614
rect 162222 464378 162306 464614
rect 162542 464378 162574 464614
rect 161954 464294 162574 464378
rect 161954 464058 161986 464294
rect 162222 464058 162306 464294
rect 162542 464058 162574 464294
rect 161954 428614 162574 464058
rect 161954 428378 161986 428614
rect 162222 428378 162306 428614
rect 162542 428378 162574 428614
rect 161954 428294 162574 428378
rect 161954 428058 161986 428294
rect 162222 428058 162306 428294
rect 162542 428058 162574 428294
rect 161954 392614 162574 428058
rect 161954 392378 161986 392614
rect 162222 392378 162306 392614
rect 162542 392378 162574 392614
rect 161954 392294 162574 392378
rect 161954 392058 161986 392294
rect 162222 392058 162306 392294
rect 162542 392058 162574 392294
rect 161954 356614 162574 392058
rect 161954 356378 161986 356614
rect 162222 356378 162306 356614
rect 162542 356378 162574 356614
rect 161954 356294 162574 356378
rect 161954 356058 161986 356294
rect 162222 356058 162306 356294
rect 162542 356058 162574 356294
rect 161954 320614 162574 356058
rect 161954 320378 161986 320614
rect 162222 320378 162306 320614
rect 162542 320378 162574 320614
rect 161954 320294 162574 320378
rect 161954 320058 161986 320294
rect 162222 320058 162306 320294
rect 162542 320058 162574 320294
rect 161954 284614 162574 320058
rect 161954 284378 161986 284614
rect 162222 284378 162306 284614
rect 162542 284378 162574 284614
rect 161954 284294 162574 284378
rect 161954 284058 161986 284294
rect 162222 284058 162306 284294
rect 162542 284058 162574 284294
rect 161954 248614 162574 284058
rect 161954 248378 161986 248614
rect 162222 248378 162306 248614
rect 162542 248378 162574 248614
rect 161954 248294 162574 248378
rect 161954 248058 161986 248294
rect 162222 248058 162306 248294
rect 162542 248058 162574 248294
rect 161954 212614 162574 248058
rect 161954 212378 161986 212614
rect 162222 212378 162306 212614
rect 162542 212378 162574 212614
rect 161954 212294 162574 212378
rect 161954 212058 161986 212294
rect 162222 212058 162306 212294
rect 162542 212058 162574 212294
rect 161954 176614 162574 212058
rect 161954 176378 161986 176614
rect 162222 176378 162306 176614
rect 162542 176378 162574 176614
rect 161954 176294 162574 176378
rect 161954 176058 161986 176294
rect 162222 176058 162306 176294
rect 162542 176058 162574 176294
rect 161954 140614 162574 176058
rect 161954 140378 161986 140614
rect 162222 140378 162306 140614
rect 162542 140378 162574 140614
rect 161954 140294 162574 140378
rect 161954 140058 161986 140294
rect 162222 140058 162306 140294
rect 162542 140058 162574 140294
rect 161954 104614 162574 140058
rect 161954 104378 161986 104614
rect 162222 104378 162306 104614
rect 162542 104378 162574 104614
rect 161954 104294 162574 104378
rect 161954 104058 161986 104294
rect 162222 104058 162306 104294
rect 162542 104058 162574 104294
rect 161954 68614 162574 104058
rect 161954 68378 161986 68614
rect 162222 68378 162306 68614
rect 162542 68378 162574 68614
rect 161954 68294 162574 68378
rect 161954 68058 161986 68294
rect 162222 68058 162306 68294
rect 162542 68058 162574 68294
rect 161954 32614 162574 68058
rect 161954 32378 161986 32614
rect 162222 32378 162306 32614
rect 162542 32378 162574 32614
rect 161954 32294 162574 32378
rect 161954 32058 161986 32294
rect 162222 32058 162306 32294
rect 162542 32058 162574 32294
rect 158234 -5382 158266 -5146
rect 158502 -5382 158586 -5146
rect 158822 -5382 158854 -5146
rect 158234 -5466 158854 -5382
rect 158234 -5702 158266 -5466
rect 158502 -5702 158586 -5466
rect 158822 -5702 158854 -5466
rect 158234 -5734 158854 -5702
rect 151954 -6342 151986 -6106
rect 152222 -6342 152306 -6106
rect 152542 -6342 152574 -6106
rect 151954 -6426 152574 -6342
rect 151954 -6662 151986 -6426
rect 152222 -6662 152306 -6426
rect 152542 -6662 152574 -6426
rect 151954 -7654 152574 -6662
rect 161954 -7066 162574 32058
rect 164514 706758 165134 707750
rect 164514 706522 164546 706758
rect 164782 706522 164866 706758
rect 165102 706522 165134 706758
rect 164514 706438 165134 706522
rect 164514 706202 164546 706438
rect 164782 706202 164866 706438
rect 165102 706202 165134 706438
rect 164514 691174 165134 706202
rect 164514 690938 164546 691174
rect 164782 690938 164866 691174
rect 165102 690938 165134 691174
rect 164514 690854 165134 690938
rect 164514 690618 164546 690854
rect 164782 690618 164866 690854
rect 165102 690618 165134 690854
rect 164514 655174 165134 690618
rect 164514 654938 164546 655174
rect 164782 654938 164866 655174
rect 165102 654938 165134 655174
rect 164514 654854 165134 654938
rect 164514 654618 164546 654854
rect 164782 654618 164866 654854
rect 165102 654618 165134 654854
rect 164514 619174 165134 654618
rect 164514 618938 164546 619174
rect 164782 618938 164866 619174
rect 165102 618938 165134 619174
rect 164514 618854 165134 618938
rect 164514 618618 164546 618854
rect 164782 618618 164866 618854
rect 165102 618618 165134 618854
rect 164514 583174 165134 618618
rect 164514 582938 164546 583174
rect 164782 582938 164866 583174
rect 165102 582938 165134 583174
rect 164514 582854 165134 582938
rect 164514 582618 164546 582854
rect 164782 582618 164866 582854
rect 165102 582618 165134 582854
rect 164514 547174 165134 582618
rect 164514 546938 164546 547174
rect 164782 546938 164866 547174
rect 165102 546938 165134 547174
rect 164514 546854 165134 546938
rect 164514 546618 164546 546854
rect 164782 546618 164866 546854
rect 165102 546618 165134 546854
rect 164514 511174 165134 546618
rect 164514 510938 164546 511174
rect 164782 510938 164866 511174
rect 165102 510938 165134 511174
rect 164514 510854 165134 510938
rect 164514 510618 164546 510854
rect 164782 510618 164866 510854
rect 165102 510618 165134 510854
rect 164514 475174 165134 510618
rect 164514 474938 164546 475174
rect 164782 474938 164866 475174
rect 165102 474938 165134 475174
rect 164514 474854 165134 474938
rect 164514 474618 164546 474854
rect 164782 474618 164866 474854
rect 165102 474618 165134 474854
rect 164514 439174 165134 474618
rect 164514 438938 164546 439174
rect 164782 438938 164866 439174
rect 165102 438938 165134 439174
rect 164514 438854 165134 438938
rect 164514 438618 164546 438854
rect 164782 438618 164866 438854
rect 165102 438618 165134 438854
rect 164514 403174 165134 438618
rect 164514 402938 164546 403174
rect 164782 402938 164866 403174
rect 165102 402938 165134 403174
rect 164514 402854 165134 402938
rect 164514 402618 164546 402854
rect 164782 402618 164866 402854
rect 165102 402618 165134 402854
rect 164514 367174 165134 402618
rect 164514 366938 164546 367174
rect 164782 366938 164866 367174
rect 165102 366938 165134 367174
rect 164514 366854 165134 366938
rect 164514 366618 164546 366854
rect 164782 366618 164866 366854
rect 165102 366618 165134 366854
rect 164514 331174 165134 366618
rect 164514 330938 164546 331174
rect 164782 330938 164866 331174
rect 165102 330938 165134 331174
rect 164514 330854 165134 330938
rect 164514 330618 164546 330854
rect 164782 330618 164866 330854
rect 165102 330618 165134 330854
rect 164514 295174 165134 330618
rect 164514 294938 164546 295174
rect 164782 294938 164866 295174
rect 165102 294938 165134 295174
rect 164514 294854 165134 294938
rect 164514 294618 164546 294854
rect 164782 294618 164866 294854
rect 165102 294618 165134 294854
rect 164514 259174 165134 294618
rect 164514 258938 164546 259174
rect 164782 258938 164866 259174
rect 165102 258938 165134 259174
rect 164514 258854 165134 258938
rect 164514 258618 164546 258854
rect 164782 258618 164866 258854
rect 165102 258618 165134 258854
rect 164514 223174 165134 258618
rect 164514 222938 164546 223174
rect 164782 222938 164866 223174
rect 165102 222938 165134 223174
rect 164514 222854 165134 222938
rect 164514 222618 164546 222854
rect 164782 222618 164866 222854
rect 165102 222618 165134 222854
rect 164514 187174 165134 222618
rect 164514 186938 164546 187174
rect 164782 186938 164866 187174
rect 165102 186938 165134 187174
rect 164514 186854 165134 186938
rect 164514 186618 164546 186854
rect 164782 186618 164866 186854
rect 165102 186618 165134 186854
rect 164514 151174 165134 186618
rect 164514 150938 164546 151174
rect 164782 150938 164866 151174
rect 165102 150938 165134 151174
rect 164514 150854 165134 150938
rect 164514 150618 164546 150854
rect 164782 150618 164866 150854
rect 165102 150618 165134 150854
rect 164514 115174 165134 150618
rect 164514 114938 164546 115174
rect 164782 114938 164866 115174
rect 165102 114938 165134 115174
rect 164514 114854 165134 114938
rect 164514 114618 164546 114854
rect 164782 114618 164866 114854
rect 165102 114618 165134 114854
rect 164514 79174 165134 114618
rect 164514 78938 164546 79174
rect 164782 78938 164866 79174
rect 165102 78938 165134 79174
rect 164514 78854 165134 78938
rect 164514 78618 164546 78854
rect 164782 78618 164866 78854
rect 165102 78618 165134 78854
rect 164514 43174 165134 78618
rect 164514 42938 164546 43174
rect 164782 42938 164866 43174
rect 165102 42938 165134 43174
rect 164514 42854 165134 42938
rect 164514 42618 164546 42854
rect 164782 42618 164866 42854
rect 165102 42618 165134 42854
rect 164514 7174 165134 42618
rect 164514 6938 164546 7174
rect 164782 6938 164866 7174
rect 165102 6938 165134 7174
rect 164514 6854 165134 6938
rect 164514 6618 164546 6854
rect 164782 6618 164866 6854
rect 165102 6618 165134 6854
rect 164514 -2266 165134 6618
rect 164514 -2502 164546 -2266
rect 164782 -2502 164866 -2266
rect 165102 -2502 165134 -2266
rect 164514 -2586 165134 -2502
rect 164514 -2822 164546 -2586
rect 164782 -2822 164866 -2586
rect 165102 -2822 165134 -2586
rect 164514 -3814 165134 -2822
rect 168234 694894 168854 708122
rect 168234 694658 168266 694894
rect 168502 694658 168586 694894
rect 168822 694658 168854 694894
rect 168234 694574 168854 694658
rect 168234 694338 168266 694574
rect 168502 694338 168586 694574
rect 168822 694338 168854 694574
rect 168234 658894 168854 694338
rect 168234 658658 168266 658894
rect 168502 658658 168586 658894
rect 168822 658658 168854 658894
rect 168234 658574 168854 658658
rect 168234 658338 168266 658574
rect 168502 658338 168586 658574
rect 168822 658338 168854 658574
rect 168234 622894 168854 658338
rect 168234 622658 168266 622894
rect 168502 622658 168586 622894
rect 168822 622658 168854 622894
rect 168234 622574 168854 622658
rect 168234 622338 168266 622574
rect 168502 622338 168586 622574
rect 168822 622338 168854 622574
rect 168234 586894 168854 622338
rect 168234 586658 168266 586894
rect 168502 586658 168586 586894
rect 168822 586658 168854 586894
rect 168234 586574 168854 586658
rect 168234 586338 168266 586574
rect 168502 586338 168586 586574
rect 168822 586338 168854 586574
rect 168234 550894 168854 586338
rect 168234 550658 168266 550894
rect 168502 550658 168586 550894
rect 168822 550658 168854 550894
rect 168234 550574 168854 550658
rect 168234 550338 168266 550574
rect 168502 550338 168586 550574
rect 168822 550338 168854 550574
rect 168234 514894 168854 550338
rect 168234 514658 168266 514894
rect 168502 514658 168586 514894
rect 168822 514658 168854 514894
rect 168234 514574 168854 514658
rect 168234 514338 168266 514574
rect 168502 514338 168586 514574
rect 168822 514338 168854 514574
rect 168234 478894 168854 514338
rect 168234 478658 168266 478894
rect 168502 478658 168586 478894
rect 168822 478658 168854 478894
rect 168234 478574 168854 478658
rect 168234 478338 168266 478574
rect 168502 478338 168586 478574
rect 168822 478338 168854 478574
rect 168234 442894 168854 478338
rect 168234 442658 168266 442894
rect 168502 442658 168586 442894
rect 168822 442658 168854 442894
rect 168234 442574 168854 442658
rect 168234 442338 168266 442574
rect 168502 442338 168586 442574
rect 168822 442338 168854 442574
rect 168234 406894 168854 442338
rect 168234 406658 168266 406894
rect 168502 406658 168586 406894
rect 168822 406658 168854 406894
rect 168234 406574 168854 406658
rect 168234 406338 168266 406574
rect 168502 406338 168586 406574
rect 168822 406338 168854 406574
rect 168234 370894 168854 406338
rect 168234 370658 168266 370894
rect 168502 370658 168586 370894
rect 168822 370658 168854 370894
rect 168234 370574 168854 370658
rect 168234 370338 168266 370574
rect 168502 370338 168586 370574
rect 168822 370338 168854 370574
rect 168234 334894 168854 370338
rect 168234 334658 168266 334894
rect 168502 334658 168586 334894
rect 168822 334658 168854 334894
rect 168234 334574 168854 334658
rect 168234 334338 168266 334574
rect 168502 334338 168586 334574
rect 168822 334338 168854 334574
rect 168234 298894 168854 334338
rect 168234 298658 168266 298894
rect 168502 298658 168586 298894
rect 168822 298658 168854 298894
rect 168234 298574 168854 298658
rect 168234 298338 168266 298574
rect 168502 298338 168586 298574
rect 168822 298338 168854 298574
rect 168234 262894 168854 298338
rect 168234 262658 168266 262894
rect 168502 262658 168586 262894
rect 168822 262658 168854 262894
rect 168234 262574 168854 262658
rect 168234 262338 168266 262574
rect 168502 262338 168586 262574
rect 168822 262338 168854 262574
rect 168234 226894 168854 262338
rect 168234 226658 168266 226894
rect 168502 226658 168586 226894
rect 168822 226658 168854 226894
rect 168234 226574 168854 226658
rect 168234 226338 168266 226574
rect 168502 226338 168586 226574
rect 168822 226338 168854 226574
rect 168234 190894 168854 226338
rect 168234 190658 168266 190894
rect 168502 190658 168586 190894
rect 168822 190658 168854 190894
rect 168234 190574 168854 190658
rect 168234 190338 168266 190574
rect 168502 190338 168586 190574
rect 168822 190338 168854 190574
rect 168234 154894 168854 190338
rect 168234 154658 168266 154894
rect 168502 154658 168586 154894
rect 168822 154658 168854 154894
rect 168234 154574 168854 154658
rect 168234 154338 168266 154574
rect 168502 154338 168586 154574
rect 168822 154338 168854 154574
rect 168234 118894 168854 154338
rect 168234 118658 168266 118894
rect 168502 118658 168586 118894
rect 168822 118658 168854 118894
rect 168234 118574 168854 118658
rect 168234 118338 168266 118574
rect 168502 118338 168586 118574
rect 168822 118338 168854 118574
rect 168234 82894 168854 118338
rect 168234 82658 168266 82894
rect 168502 82658 168586 82894
rect 168822 82658 168854 82894
rect 168234 82574 168854 82658
rect 168234 82338 168266 82574
rect 168502 82338 168586 82574
rect 168822 82338 168854 82574
rect 168234 46894 168854 82338
rect 168234 46658 168266 46894
rect 168502 46658 168586 46894
rect 168822 46658 168854 46894
rect 168234 46574 168854 46658
rect 168234 46338 168266 46574
rect 168502 46338 168586 46574
rect 168822 46338 168854 46574
rect 168234 10894 168854 46338
rect 168234 10658 168266 10894
rect 168502 10658 168586 10894
rect 168822 10658 168854 10894
rect 168234 10574 168854 10658
rect 168234 10338 168266 10574
rect 168502 10338 168586 10574
rect 168822 10338 168854 10574
rect 168234 -4186 168854 10338
rect 170794 705798 171414 705830
rect 170794 705562 170826 705798
rect 171062 705562 171146 705798
rect 171382 705562 171414 705798
rect 170794 705478 171414 705562
rect 170794 705242 170826 705478
rect 171062 705242 171146 705478
rect 171382 705242 171414 705478
rect 170794 669454 171414 705242
rect 170794 669218 170826 669454
rect 171062 669218 171146 669454
rect 171382 669218 171414 669454
rect 170794 669134 171414 669218
rect 170794 668898 170826 669134
rect 171062 668898 171146 669134
rect 171382 668898 171414 669134
rect 170794 633454 171414 668898
rect 170794 633218 170826 633454
rect 171062 633218 171146 633454
rect 171382 633218 171414 633454
rect 170794 633134 171414 633218
rect 170794 632898 170826 633134
rect 171062 632898 171146 633134
rect 171382 632898 171414 633134
rect 170794 597454 171414 632898
rect 170794 597218 170826 597454
rect 171062 597218 171146 597454
rect 171382 597218 171414 597454
rect 170794 597134 171414 597218
rect 170794 596898 170826 597134
rect 171062 596898 171146 597134
rect 171382 596898 171414 597134
rect 170794 561454 171414 596898
rect 170794 561218 170826 561454
rect 171062 561218 171146 561454
rect 171382 561218 171414 561454
rect 170794 561134 171414 561218
rect 170794 560898 170826 561134
rect 171062 560898 171146 561134
rect 171382 560898 171414 561134
rect 170794 525454 171414 560898
rect 170794 525218 170826 525454
rect 171062 525218 171146 525454
rect 171382 525218 171414 525454
rect 170794 525134 171414 525218
rect 170794 524898 170826 525134
rect 171062 524898 171146 525134
rect 171382 524898 171414 525134
rect 170794 489454 171414 524898
rect 170794 489218 170826 489454
rect 171062 489218 171146 489454
rect 171382 489218 171414 489454
rect 170794 489134 171414 489218
rect 170794 488898 170826 489134
rect 171062 488898 171146 489134
rect 171382 488898 171414 489134
rect 170794 453454 171414 488898
rect 170794 453218 170826 453454
rect 171062 453218 171146 453454
rect 171382 453218 171414 453454
rect 170794 453134 171414 453218
rect 170794 452898 170826 453134
rect 171062 452898 171146 453134
rect 171382 452898 171414 453134
rect 170794 417454 171414 452898
rect 170794 417218 170826 417454
rect 171062 417218 171146 417454
rect 171382 417218 171414 417454
rect 170794 417134 171414 417218
rect 170794 416898 170826 417134
rect 171062 416898 171146 417134
rect 171382 416898 171414 417134
rect 170794 381454 171414 416898
rect 170794 381218 170826 381454
rect 171062 381218 171146 381454
rect 171382 381218 171414 381454
rect 170794 381134 171414 381218
rect 170794 380898 170826 381134
rect 171062 380898 171146 381134
rect 171382 380898 171414 381134
rect 170794 345454 171414 380898
rect 170794 345218 170826 345454
rect 171062 345218 171146 345454
rect 171382 345218 171414 345454
rect 170794 345134 171414 345218
rect 170794 344898 170826 345134
rect 171062 344898 171146 345134
rect 171382 344898 171414 345134
rect 170794 309454 171414 344898
rect 170794 309218 170826 309454
rect 171062 309218 171146 309454
rect 171382 309218 171414 309454
rect 170794 309134 171414 309218
rect 170794 308898 170826 309134
rect 171062 308898 171146 309134
rect 171382 308898 171414 309134
rect 170794 273454 171414 308898
rect 170794 273218 170826 273454
rect 171062 273218 171146 273454
rect 171382 273218 171414 273454
rect 170794 273134 171414 273218
rect 170794 272898 170826 273134
rect 171062 272898 171146 273134
rect 171382 272898 171414 273134
rect 170794 237454 171414 272898
rect 170794 237218 170826 237454
rect 171062 237218 171146 237454
rect 171382 237218 171414 237454
rect 170794 237134 171414 237218
rect 170794 236898 170826 237134
rect 171062 236898 171146 237134
rect 171382 236898 171414 237134
rect 170794 201454 171414 236898
rect 170794 201218 170826 201454
rect 171062 201218 171146 201454
rect 171382 201218 171414 201454
rect 170794 201134 171414 201218
rect 170794 200898 170826 201134
rect 171062 200898 171146 201134
rect 171382 200898 171414 201134
rect 170794 165454 171414 200898
rect 170794 165218 170826 165454
rect 171062 165218 171146 165454
rect 171382 165218 171414 165454
rect 170794 165134 171414 165218
rect 170794 164898 170826 165134
rect 171062 164898 171146 165134
rect 171382 164898 171414 165134
rect 170794 129454 171414 164898
rect 170794 129218 170826 129454
rect 171062 129218 171146 129454
rect 171382 129218 171414 129454
rect 170794 129134 171414 129218
rect 170794 128898 170826 129134
rect 171062 128898 171146 129134
rect 171382 128898 171414 129134
rect 170794 93454 171414 128898
rect 170794 93218 170826 93454
rect 171062 93218 171146 93454
rect 171382 93218 171414 93454
rect 170794 93134 171414 93218
rect 170794 92898 170826 93134
rect 171062 92898 171146 93134
rect 171382 92898 171414 93134
rect 170794 57454 171414 92898
rect 170794 57218 170826 57454
rect 171062 57218 171146 57454
rect 171382 57218 171414 57454
rect 170794 57134 171414 57218
rect 170794 56898 170826 57134
rect 171062 56898 171146 57134
rect 171382 56898 171414 57134
rect 170794 21454 171414 56898
rect 170794 21218 170826 21454
rect 171062 21218 171146 21454
rect 171382 21218 171414 21454
rect 170794 21134 171414 21218
rect 170794 20898 170826 21134
rect 171062 20898 171146 21134
rect 171382 20898 171414 21134
rect 170794 -1306 171414 20898
rect 170794 -1542 170826 -1306
rect 171062 -1542 171146 -1306
rect 171382 -1542 171414 -1306
rect 170794 -1626 171414 -1542
rect 170794 -1862 170826 -1626
rect 171062 -1862 171146 -1626
rect 171382 -1862 171414 -1626
rect 170794 -1894 171414 -1862
rect 171954 698614 172574 710042
rect 181954 711558 182574 711590
rect 181954 711322 181986 711558
rect 182222 711322 182306 711558
rect 182542 711322 182574 711558
rect 181954 711238 182574 711322
rect 181954 711002 181986 711238
rect 182222 711002 182306 711238
rect 182542 711002 182574 711238
rect 178234 709638 178854 709670
rect 178234 709402 178266 709638
rect 178502 709402 178586 709638
rect 178822 709402 178854 709638
rect 178234 709318 178854 709402
rect 178234 709082 178266 709318
rect 178502 709082 178586 709318
rect 178822 709082 178854 709318
rect 171954 698378 171986 698614
rect 172222 698378 172306 698614
rect 172542 698378 172574 698614
rect 171954 698294 172574 698378
rect 171954 698058 171986 698294
rect 172222 698058 172306 698294
rect 172542 698058 172574 698294
rect 171954 662614 172574 698058
rect 171954 662378 171986 662614
rect 172222 662378 172306 662614
rect 172542 662378 172574 662614
rect 171954 662294 172574 662378
rect 171954 662058 171986 662294
rect 172222 662058 172306 662294
rect 172542 662058 172574 662294
rect 171954 626614 172574 662058
rect 171954 626378 171986 626614
rect 172222 626378 172306 626614
rect 172542 626378 172574 626614
rect 171954 626294 172574 626378
rect 171954 626058 171986 626294
rect 172222 626058 172306 626294
rect 172542 626058 172574 626294
rect 171954 590614 172574 626058
rect 171954 590378 171986 590614
rect 172222 590378 172306 590614
rect 172542 590378 172574 590614
rect 171954 590294 172574 590378
rect 171954 590058 171986 590294
rect 172222 590058 172306 590294
rect 172542 590058 172574 590294
rect 171954 554614 172574 590058
rect 171954 554378 171986 554614
rect 172222 554378 172306 554614
rect 172542 554378 172574 554614
rect 171954 554294 172574 554378
rect 171954 554058 171986 554294
rect 172222 554058 172306 554294
rect 172542 554058 172574 554294
rect 171954 518614 172574 554058
rect 171954 518378 171986 518614
rect 172222 518378 172306 518614
rect 172542 518378 172574 518614
rect 171954 518294 172574 518378
rect 171954 518058 171986 518294
rect 172222 518058 172306 518294
rect 172542 518058 172574 518294
rect 171954 482614 172574 518058
rect 171954 482378 171986 482614
rect 172222 482378 172306 482614
rect 172542 482378 172574 482614
rect 171954 482294 172574 482378
rect 171954 482058 171986 482294
rect 172222 482058 172306 482294
rect 172542 482058 172574 482294
rect 171954 446614 172574 482058
rect 171954 446378 171986 446614
rect 172222 446378 172306 446614
rect 172542 446378 172574 446614
rect 171954 446294 172574 446378
rect 171954 446058 171986 446294
rect 172222 446058 172306 446294
rect 172542 446058 172574 446294
rect 171954 410614 172574 446058
rect 171954 410378 171986 410614
rect 172222 410378 172306 410614
rect 172542 410378 172574 410614
rect 171954 410294 172574 410378
rect 171954 410058 171986 410294
rect 172222 410058 172306 410294
rect 172542 410058 172574 410294
rect 171954 374614 172574 410058
rect 171954 374378 171986 374614
rect 172222 374378 172306 374614
rect 172542 374378 172574 374614
rect 171954 374294 172574 374378
rect 171954 374058 171986 374294
rect 172222 374058 172306 374294
rect 172542 374058 172574 374294
rect 171954 338614 172574 374058
rect 171954 338378 171986 338614
rect 172222 338378 172306 338614
rect 172542 338378 172574 338614
rect 171954 338294 172574 338378
rect 171954 338058 171986 338294
rect 172222 338058 172306 338294
rect 172542 338058 172574 338294
rect 171954 302614 172574 338058
rect 171954 302378 171986 302614
rect 172222 302378 172306 302614
rect 172542 302378 172574 302614
rect 171954 302294 172574 302378
rect 171954 302058 171986 302294
rect 172222 302058 172306 302294
rect 172542 302058 172574 302294
rect 171954 266614 172574 302058
rect 171954 266378 171986 266614
rect 172222 266378 172306 266614
rect 172542 266378 172574 266614
rect 171954 266294 172574 266378
rect 171954 266058 171986 266294
rect 172222 266058 172306 266294
rect 172542 266058 172574 266294
rect 171954 230614 172574 266058
rect 171954 230378 171986 230614
rect 172222 230378 172306 230614
rect 172542 230378 172574 230614
rect 171954 230294 172574 230378
rect 171954 230058 171986 230294
rect 172222 230058 172306 230294
rect 172542 230058 172574 230294
rect 171954 194614 172574 230058
rect 171954 194378 171986 194614
rect 172222 194378 172306 194614
rect 172542 194378 172574 194614
rect 171954 194294 172574 194378
rect 171954 194058 171986 194294
rect 172222 194058 172306 194294
rect 172542 194058 172574 194294
rect 171954 158614 172574 194058
rect 171954 158378 171986 158614
rect 172222 158378 172306 158614
rect 172542 158378 172574 158614
rect 171954 158294 172574 158378
rect 171954 158058 171986 158294
rect 172222 158058 172306 158294
rect 172542 158058 172574 158294
rect 171954 122614 172574 158058
rect 171954 122378 171986 122614
rect 172222 122378 172306 122614
rect 172542 122378 172574 122614
rect 171954 122294 172574 122378
rect 171954 122058 171986 122294
rect 172222 122058 172306 122294
rect 172542 122058 172574 122294
rect 171954 86614 172574 122058
rect 171954 86378 171986 86614
rect 172222 86378 172306 86614
rect 172542 86378 172574 86614
rect 171954 86294 172574 86378
rect 171954 86058 171986 86294
rect 172222 86058 172306 86294
rect 172542 86058 172574 86294
rect 171954 50614 172574 86058
rect 171954 50378 171986 50614
rect 172222 50378 172306 50614
rect 172542 50378 172574 50614
rect 171954 50294 172574 50378
rect 171954 50058 171986 50294
rect 172222 50058 172306 50294
rect 172542 50058 172574 50294
rect 171954 14614 172574 50058
rect 171954 14378 171986 14614
rect 172222 14378 172306 14614
rect 172542 14378 172574 14614
rect 171954 14294 172574 14378
rect 171954 14058 171986 14294
rect 172222 14058 172306 14294
rect 172542 14058 172574 14294
rect 168234 -4422 168266 -4186
rect 168502 -4422 168586 -4186
rect 168822 -4422 168854 -4186
rect 168234 -4506 168854 -4422
rect 168234 -4742 168266 -4506
rect 168502 -4742 168586 -4506
rect 168822 -4742 168854 -4506
rect 168234 -5734 168854 -4742
rect 161954 -7302 161986 -7066
rect 162222 -7302 162306 -7066
rect 162542 -7302 162574 -7066
rect 161954 -7386 162574 -7302
rect 161954 -7622 161986 -7386
rect 162222 -7622 162306 -7386
rect 162542 -7622 162574 -7386
rect 161954 -7654 162574 -7622
rect 171954 -6106 172574 14058
rect 174514 707718 175134 707750
rect 174514 707482 174546 707718
rect 174782 707482 174866 707718
rect 175102 707482 175134 707718
rect 174514 707398 175134 707482
rect 174514 707162 174546 707398
rect 174782 707162 174866 707398
rect 175102 707162 175134 707398
rect 174514 673174 175134 707162
rect 174514 672938 174546 673174
rect 174782 672938 174866 673174
rect 175102 672938 175134 673174
rect 174514 672854 175134 672938
rect 174514 672618 174546 672854
rect 174782 672618 174866 672854
rect 175102 672618 175134 672854
rect 174514 637174 175134 672618
rect 174514 636938 174546 637174
rect 174782 636938 174866 637174
rect 175102 636938 175134 637174
rect 174514 636854 175134 636938
rect 174514 636618 174546 636854
rect 174782 636618 174866 636854
rect 175102 636618 175134 636854
rect 174514 601174 175134 636618
rect 174514 600938 174546 601174
rect 174782 600938 174866 601174
rect 175102 600938 175134 601174
rect 174514 600854 175134 600938
rect 174514 600618 174546 600854
rect 174782 600618 174866 600854
rect 175102 600618 175134 600854
rect 174514 565174 175134 600618
rect 174514 564938 174546 565174
rect 174782 564938 174866 565174
rect 175102 564938 175134 565174
rect 174514 564854 175134 564938
rect 174514 564618 174546 564854
rect 174782 564618 174866 564854
rect 175102 564618 175134 564854
rect 174514 529174 175134 564618
rect 174514 528938 174546 529174
rect 174782 528938 174866 529174
rect 175102 528938 175134 529174
rect 174514 528854 175134 528938
rect 174514 528618 174546 528854
rect 174782 528618 174866 528854
rect 175102 528618 175134 528854
rect 174514 493174 175134 528618
rect 174514 492938 174546 493174
rect 174782 492938 174866 493174
rect 175102 492938 175134 493174
rect 174514 492854 175134 492938
rect 174514 492618 174546 492854
rect 174782 492618 174866 492854
rect 175102 492618 175134 492854
rect 174514 457174 175134 492618
rect 174514 456938 174546 457174
rect 174782 456938 174866 457174
rect 175102 456938 175134 457174
rect 174514 456854 175134 456938
rect 174514 456618 174546 456854
rect 174782 456618 174866 456854
rect 175102 456618 175134 456854
rect 174514 421174 175134 456618
rect 174514 420938 174546 421174
rect 174782 420938 174866 421174
rect 175102 420938 175134 421174
rect 174514 420854 175134 420938
rect 174514 420618 174546 420854
rect 174782 420618 174866 420854
rect 175102 420618 175134 420854
rect 174514 385174 175134 420618
rect 174514 384938 174546 385174
rect 174782 384938 174866 385174
rect 175102 384938 175134 385174
rect 174514 384854 175134 384938
rect 174514 384618 174546 384854
rect 174782 384618 174866 384854
rect 175102 384618 175134 384854
rect 174514 349174 175134 384618
rect 174514 348938 174546 349174
rect 174782 348938 174866 349174
rect 175102 348938 175134 349174
rect 174514 348854 175134 348938
rect 174514 348618 174546 348854
rect 174782 348618 174866 348854
rect 175102 348618 175134 348854
rect 174514 313174 175134 348618
rect 174514 312938 174546 313174
rect 174782 312938 174866 313174
rect 175102 312938 175134 313174
rect 174514 312854 175134 312938
rect 174514 312618 174546 312854
rect 174782 312618 174866 312854
rect 175102 312618 175134 312854
rect 174514 277174 175134 312618
rect 174514 276938 174546 277174
rect 174782 276938 174866 277174
rect 175102 276938 175134 277174
rect 174514 276854 175134 276938
rect 174514 276618 174546 276854
rect 174782 276618 174866 276854
rect 175102 276618 175134 276854
rect 174514 241174 175134 276618
rect 174514 240938 174546 241174
rect 174782 240938 174866 241174
rect 175102 240938 175134 241174
rect 174514 240854 175134 240938
rect 174514 240618 174546 240854
rect 174782 240618 174866 240854
rect 175102 240618 175134 240854
rect 174514 205174 175134 240618
rect 174514 204938 174546 205174
rect 174782 204938 174866 205174
rect 175102 204938 175134 205174
rect 174514 204854 175134 204938
rect 174514 204618 174546 204854
rect 174782 204618 174866 204854
rect 175102 204618 175134 204854
rect 174514 169174 175134 204618
rect 174514 168938 174546 169174
rect 174782 168938 174866 169174
rect 175102 168938 175134 169174
rect 174514 168854 175134 168938
rect 174514 168618 174546 168854
rect 174782 168618 174866 168854
rect 175102 168618 175134 168854
rect 174514 133174 175134 168618
rect 174514 132938 174546 133174
rect 174782 132938 174866 133174
rect 175102 132938 175134 133174
rect 174514 132854 175134 132938
rect 174514 132618 174546 132854
rect 174782 132618 174866 132854
rect 175102 132618 175134 132854
rect 174514 97174 175134 132618
rect 174514 96938 174546 97174
rect 174782 96938 174866 97174
rect 175102 96938 175134 97174
rect 174514 96854 175134 96938
rect 174514 96618 174546 96854
rect 174782 96618 174866 96854
rect 175102 96618 175134 96854
rect 174514 61174 175134 96618
rect 174514 60938 174546 61174
rect 174782 60938 174866 61174
rect 175102 60938 175134 61174
rect 174514 60854 175134 60938
rect 174514 60618 174546 60854
rect 174782 60618 174866 60854
rect 175102 60618 175134 60854
rect 174514 25174 175134 60618
rect 174514 24938 174546 25174
rect 174782 24938 174866 25174
rect 175102 24938 175134 25174
rect 174514 24854 175134 24938
rect 174514 24618 174546 24854
rect 174782 24618 174866 24854
rect 175102 24618 175134 24854
rect 174514 -3226 175134 24618
rect 174514 -3462 174546 -3226
rect 174782 -3462 174866 -3226
rect 175102 -3462 175134 -3226
rect 174514 -3546 175134 -3462
rect 174514 -3782 174546 -3546
rect 174782 -3782 174866 -3546
rect 175102 -3782 175134 -3546
rect 174514 -3814 175134 -3782
rect 178234 676894 178854 709082
rect 178234 676658 178266 676894
rect 178502 676658 178586 676894
rect 178822 676658 178854 676894
rect 178234 676574 178854 676658
rect 178234 676338 178266 676574
rect 178502 676338 178586 676574
rect 178822 676338 178854 676574
rect 178234 640894 178854 676338
rect 178234 640658 178266 640894
rect 178502 640658 178586 640894
rect 178822 640658 178854 640894
rect 178234 640574 178854 640658
rect 178234 640338 178266 640574
rect 178502 640338 178586 640574
rect 178822 640338 178854 640574
rect 178234 604894 178854 640338
rect 178234 604658 178266 604894
rect 178502 604658 178586 604894
rect 178822 604658 178854 604894
rect 178234 604574 178854 604658
rect 178234 604338 178266 604574
rect 178502 604338 178586 604574
rect 178822 604338 178854 604574
rect 178234 568894 178854 604338
rect 178234 568658 178266 568894
rect 178502 568658 178586 568894
rect 178822 568658 178854 568894
rect 178234 568574 178854 568658
rect 178234 568338 178266 568574
rect 178502 568338 178586 568574
rect 178822 568338 178854 568574
rect 178234 532894 178854 568338
rect 178234 532658 178266 532894
rect 178502 532658 178586 532894
rect 178822 532658 178854 532894
rect 178234 532574 178854 532658
rect 178234 532338 178266 532574
rect 178502 532338 178586 532574
rect 178822 532338 178854 532574
rect 178234 496894 178854 532338
rect 178234 496658 178266 496894
rect 178502 496658 178586 496894
rect 178822 496658 178854 496894
rect 178234 496574 178854 496658
rect 178234 496338 178266 496574
rect 178502 496338 178586 496574
rect 178822 496338 178854 496574
rect 178234 460894 178854 496338
rect 178234 460658 178266 460894
rect 178502 460658 178586 460894
rect 178822 460658 178854 460894
rect 178234 460574 178854 460658
rect 178234 460338 178266 460574
rect 178502 460338 178586 460574
rect 178822 460338 178854 460574
rect 178234 424894 178854 460338
rect 178234 424658 178266 424894
rect 178502 424658 178586 424894
rect 178822 424658 178854 424894
rect 178234 424574 178854 424658
rect 178234 424338 178266 424574
rect 178502 424338 178586 424574
rect 178822 424338 178854 424574
rect 178234 388894 178854 424338
rect 178234 388658 178266 388894
rect 178502 388658 178586 388894
rect 178822 388658 178854 388894
rect 178234 388574 178854 388658
rect 178234 388338 178266 388574
rect 178502 388338 178586 388574
rect 178822 388338 178854 388574
rect 178234 352894 178854 388338
rect 178234 352658 178266 352894
rect 178502 352658 178586 352894
rect 178822 352658 178854 352894
rect 178234 352574 178854 352658
rect 178234 352338 178266 352574
rect 178502 352338 178586 352574
rect 178822 352338 178854 352574
rect 178234 316894 178854 352338
rect 178234 316658 178266 316894
rect 178502 316658 178586 316894
rect 178822 316658 178854 316894
rect 178234 316574 178854 316658
rect 178234 316338 178266 316574
rect 178502 316338 178586 316574
rect 178822 316338 178854 316574
rect 178234 280894 178854 316338
rect 178234 280658 178266 280894
rect 178502 280658 178586 280894
rect 178822 280658 178854 280894
rect 178234 280574 178854 280658
rect 178234 280338 178266 280574
rect 178502 280338 178586 280574
rect 178822 280338 178854 280574
rect 178234 244894 178854 280338
rect 178234 244658 178266 244894
rect 178502 244658 178586 244894
rect 178822 244658 178854 244894
rect 178234 244574 178854 244658
rect 178234 244338 178266 244574
rect 178502 244338 178586 244574
rect 178822 244338 178854 244574
rect 178234 208894 178854 244338
rect 178234 208658 178266 208894
rect 178502 208658 178586 208894
rect 178822 208658 178854 208894
rect 178234 208574 178854 208658
rect 178234 208338 178266 208574
rect 178502 208338 178586 208574
rect 178822 208338 178854 208574
rect 178234 172894 178854 208338
rect 178234 172658 178266 172894
rect 178502 172658 178586 172894
rect 178822 172658 178854 172894
rect 178234 172574 178854 172658
rect 178234 172338 178266 172574
rect 178502 172338 178586 172574
rect 178822 172338 178854 172574
rect 178234 136894 178854 172338
rect 178234 136658 178266 136894
rect 178502 136658 178586 136894
rect 178822 136658 178854 136894
rect 178234 136574 178854 136658
rect 178234 136338 178266 136574
rect 178502 136338 178586 136574
rect 178822 136338 178854 136574
rect 178234 100894 178854 136338
rect 178234 100658 178266 100894
rect 178502 100658 178586 100894
rect 178822 100658 178854 100894
rect 178234 100574 178854 100658
rect 178234 100338 178266 100574
rect 178502 100338 178586 100574
rect 178822 100338 178854 100574
rect 178234 64894 178854 100338
rect 178234 64658 178266 64894
rect 178502 64658 178586 64894
rect 178822 64658 178854 64894
rect 178234 64574 178854 64658
rect 178234 64338 178266 64574
rect 178502 64338 178586 64574
rect 178822 64338 178854 64574
rect 178234 28894 178854 64338
rect 178234 28658 178266 28894
rect 178502 28658 178586 28894
rect 178822 28658 178854 28894
rect 178234 28574 178854 28658
rect 178234 28338 178266 28574
rect 178502 28338 178586 28574
rect 178822 28338 178854 28574
rect 178234 -5146 178854 28338
rect 180794 704838 181414 705830
rect 180794 704602 180826 704838
rect 181062 704602 181146 704838
rect 181382 704602 181414 704838
rect 180794 704518 181414 704602
rect 180794 704282 180826 704518
rect 181062 704282 181146 704518
rect 181382 704282 181414 704518
rect 180794 687454 181414 704282
rect 180794 687218 180826 687454
rect 181062 687218 181146 687454
rect 181382 687218 181414 687454
rect 180794 687134 181414 687218
rect 180794 686898 180826 687134
rect 181062 686898 181146 687134
rect 181382 686898 181414 687134
rect 180794 651454 181414 686898
rect 180794 651218 180826 651454
rect 181062 651218 181146 651454
rect 181382 651218 181414 651454
rect 180794 651134 181414 651218
rect 180794 650898 180826 651134
rect 181062 650898 181146 651134
rect 181382 650898 181414 651134
rect 180794 615454 181414 650898
rect 180794 615218 180826 615454
rect 181062 615218 181146 615454
rect 181382 615218 181414 615454
rect 180794 615134 181414 615218
rect 180794 614898 180826 615134
rect 181062 614898 181146 615134
rect 181382 614898 181414 615134
rect 180794 579454 181414 614898
rect 180794 579218 180826 579454
rect 181062 579218 181146 579454
rect 181382 579218 181414 579454
rect 180794 579134 181414 579218
rect 180794 578898 180826 579134
rect 181062 578898 181146 579134
rect 181382 578898 181414 579134
rect 180794 543454 181414 578898
rect 180794 543218 180826 543454
rect 181062 543218 181146 543454
rect 181382 543218 181414 543454
rect 180794 543134 181414 543218
rect 180794 542898 180826 543134
rect 181062 542898 181146 543134
rect 181382 542898 181414 543134
rect 180794 507454 181414 542898
rect 180794 507218 180826 507454
rect 181062 507218 181146 507454
rect 181382 507218 181414 507454
rect 180794 507134 181414 507218
rect 180794 506898 180826 507134
rect 181062 506898 181146 507134
rect 181382 506898 181414 507134
rect 180794 471454 181414 506898
rect 180794 471218 180826 471454
rect 181062 471218 181146 471454
rect 181382 471218 181414 471454
rect 180794 471134 181414 471218
rect 180794 470898 180826 471134
rect 181062 470898 181146 471134
rect 181382 470898 181414 471134
rect 180794 435454 181414 470898
rect 180794 435218 180826 435454
rect 181062 435218 181146 435454
rect 181382 435218 181414 435454
rect 180794 435134 181414 435218
rect 180794 434898 180826 435134
rect 181062 434898 181146 435134
rect 181382 434898 181414 435134
rect 180794 399454 181414 434898
rect 180794 399218 180826 399454
rect 181062 399218 181146 399454
rect 181382 399218 181414 399454
rect 180794 399134 181414 399218
rect 180794 398898 180826 399134
rect 181062 398898 181146 399134
rect 181382 398898 181414 399134
rect 180794 363454 181414 398898
rect 180794 363218 180826 363454
rect 181062 363218 181146 363454
rect 181382 363218 181414 363454
rect 180794 363134 181414 363218
rect 180794 362898 180826 363134
rect 181062 362898 181146 363134
rect 181382 362898 181414 363134
rect 180794 327454 181414 362898
rect 180794 327218 180826 327454
rect 181062 327218 181146 327454
rect 181382 327218 181414 327454
rect 180794 327134 181414 327218
rect 180794 326898 180826 327134
rect 181062 326898 181146 327134
rect 181382 326898 181414 327134
rect 180794 291454 181414 326898
rect 180794 291218 180826 291454
rect 181062 291218 181146 291454
rect 181382 291218 181414 291454
rect 180794 291134 181414 291218
rect 180794 290898 180826 291134
rect 181062 290898 181146 291134
rect 181382 290898 181414 291134
rect 180794 255454 181414 290898
rect 180794 255218 180826 255454
rect 181062 255218 181146 255454
rect 181382 255218 181414 255454
rect 180794 255134 181414 255218
rect 180794 254898 180826 255134
rect 181062 254898 181146 255134
rect 181382 254898 181414 255134
rect 180794 219454 181414 254898
rect 180794 219218 180826 219454
rect 181062 219218 181146 219454
rect 181382 219218 181414 219454
rect 180794 219134 181414 219218
rect 180794 218898 180826 219134
rect 181062 218898 181146 219134
rect 181382 218898 181414 219134
rect 180794 183454 181414 218898
rect 180794 183218 180826 183454
rect 181062 183218 181146 183454
rect 181382 183218 181414 183454
rect 180794 183134 181414 183218
rect 180794 182898 180826 183134
rect 181062 182898 181146 183134
rect 181382 182898 181414 183134
rect 180794 147454 181414 182898
rect 180794 147218 180826 147454
rect 181062 147218 181146 147454
rect 181382 147218 181414 147454
rect 180794 147134 181414 147218
rect 180794 146898 180826 147134
rect 181062 146898 181146 147134
rect 181382 146898 181414 147134
rect 180794 111454 181414 146898
rect 180794 111218 180826 111454
rect 181062 111218 181146 111454
rect 181382 111218 181414 111454
rect 180794 111134 181414 111218
rect 180794 110898 180826 111134
rect 181062 110898 181146 111134
rect 181382 110898 181414 111134
rect 180794 75454 181414 110898
rect 180794 75218 180826 75454
rect 181062 75218 181146 75454
rect 181382 75218 181414 75454
rect 180794 75134 181414 75218
rect 180794 74898 180826 75134
rect 181062 74898 181146 75134
rect 181382 74898 181414 75134
rect 180794 39454 181414 74898
rect 180794 39218 180826 39454
rect 181062 39218 181146 39454
rect 181382 39218 181414 39454
rect 180794 39134 181414 39218
rect 180794 38898 180826 39134
rect 181062 38898 181146 39134
rect 181382 38898 181414 39134
rect 180794 3454 181414 38898
rect 180794 3218 180826 3454
rect 181062 3218 181146 3454
rect 181382 3218 181414 3454
rect 180794 3134 181414 3218
rect 180794 2898 180826 3134
rect 181062 2898 181146 3134
rect 181382 2898 181414 3134
rect 180794 -346 181414 2898
rect 180794 -582 180826 -346
rect 181062 -582 181146 -346
rect 181382 -582 181414 -346
rect 180794 -666 181414 -582
rect 180794 -902 180826 -666
rect 181062 -902 181146 -666
rect 181382 -902 181414 -666
rect 180794 -1894 181414 -902
rect 181954 680614 182574 711002
rect 191954 710598 192574 711590
rect 191954 710362 191986 710598
rect 192222 710362 192306 710598
rect 192542 710362 192574 710598
rect 191954 710278 192574 710362
rect 191954 710042 191986 710278
rect 192222 710042 192306 710278
rect 192542 710042 192574 710278
rect 188234 708678 188854 709670
rect 188234 708442 188266 708678
rect 188502 708442 188586 708678
rect 188822 708442 188854 708678
rect 188234 708358 188854 708442
rect 188234 708122 188266 708358
rect 188502 708122 188586 708358
rect 188822 708122 188854 708358
rect 181954 680378 181986 680614
rect 182222 680378 182306 680614
rect 182542 680378 182574 680614
rect 181954 680294 182574 680378
rect 181954 680058 181986 680294
rect 182222 680058 182306 680294
rect 182542 680058 182574 680294
rect 181954 644614 182574 680058
rect 181954 644378 181986 644614
rect 182222 644378 182306 644614
rect 182542 644378 182574 644614
rect 181954 644294 182574 644378
rect 181954 644058 181986 644294
rect 182222 644058 182306 644294
rect 182542 644058 182574 644294
rect 181954 608614 182574 644058
rect 181954 608378 181986 608614
rect 182222 608378 182306 608614
rect 182542 608378 182574 608614
rect 181954 608294 182574 608378
rect 181954 608058 181986 608294
rect 182222 608058 182306 608294
rect 182542 608058 182574 608294
rect 181954 572614 182574 608058
rect 181954 572378 181986 572614
rect 182222 572378 182306 572614
rect 182542 572378 182574 572614
rect 181954 572294 182574 572378
rect 181954 572058 181986 572294
rect 182222 572058 182306 572294
rect 182542 572058 182574 572294
rect 181954 536614 182574 572058
rect 181954 536378 181986 536614
rect 182222 536378 182306 536614
rect 182542 536378 182574 536614
rect 181954 536294 182574 536378
rect 181954 536058 181986 536294
rect 182222 536058 182306 536294
rect 182542 536058 182574 536294
rect 181954 500614 182574 536058
rect 181954 500378 181986 500614
rect 182222 500378 182306 500614
rect 182542 500378 182574 500614
rect 181954 500294 182574 500378
rect 181954 500058 181986 500294
rect 182222 500058 182306 500294
rect 182542 500058 182574 500294
rect 181954 464614 182574 500058
rect 181954 464378 181986 464614
rect 182222 464378 182306 464614
rect 182542 464378 182574 464614
rect 181954 464294 182574 464378
rect 181954 464058 181986 464294
rect 182222 464058 182306 464294
rect 182542 464058 182574 464294
rect 181954 428614 182574 464058
rect 181954 428378 181986 428614
rect 182222 428378 182306 428614
rect 182542 428378 182574 428614
rect 181954 428294 182574 428378
rect 181954 428058 181986 428294
rect 182222 428058 182306 428294
rect 182542 428058 182574 428294
rect 181954 392614 182574 428058
rect 181954 392378 181986 392614
rect 182222 392378 182306 392614
rect 182542 392378 182574 392614
rect 181954 392294 182574 392378
rect 181954 392058 181986 392294
rect 182222 392058 182306 392294
rect 182542 392058 182574 392294
rect 181954 356614 182574 392058
rect 181954 356378 181986 356614
rect 182222 356378 182306 356614
rect 182542 356378 182574 356614
rect 181954 356294 182574 356378
rect 181954 356058 181986 356294
rect 182222 356058 182306 356294
rect 182542 356058 182574 356294
rect 181954 320614 182574 356058
rect 181954 320378 181986 320614
rect 182222 320378 182306 320614
rect 182542 320378 182574 320614
rect 181954 320294 182574 320378
rect 181954 320058 181986 320294
rect 182222 320058 182306 320294
rect 182542 320058 182574 320294
rect 181954 284614 182574 320058
rect 181954 284378 181986 284614
rect 182222 284378 182306 284614
rect 182542 284378 182574 284614
rect 181954 284294 182574 284378
rect 181954 284058 181986 284294
rect 182222 284058 182306 284294
rect 182542 284058 182574 284294
rect 181954 248614 182574 284058
rect 181954 248378 181986 248614
rect 182222 248378 182306 248614
rect 182542 248378 182574 248614
rect 181954 248294 182574 248378
rect 181954 248058 181986 248294
rect 182222 248058 182306 248294
rect 182542 248058 182574 248294
rect 181954 212614 182574 248058
rect 181954 212378 181986 212614
rect 182222 212378 182306 212614
rect 182542 212378 182574 212614
rect 181954 212294 182574 212378
rect 181954 212058 181986 212294
rect 182222 212058 182306 212294
rect 182542 212058 182574 212294
rect 181954 176614 182574 212058
rect 181954 176378 181986 176614
rect 182222 176378 182306 176614
rect 182542 176378 182574 176614
rect 181954 176294 182574 176378
rect 181954 176058 181986 176294
rect 182222 176058 182306 176294
rect 182542 176058 182574 176294
rect 181954 140614 182574 176058
rect 181954 140378 181986 140614
rect 182222 140378 182306 140614
rect 182542 140378 182574 140614
rect 181954 140294 182574 140378
rect 181954 140058 181986 140294
rect 182222 140058 182306 140294
rect 182542 140058 182574 140294
rect 181954 104614 182574 140058
rect 181954 104378 181986 104614
rect 182222 104378 182306 104614
rect 182542 104378 182574 104614
rect 181954 104294 182574 104378
rect 181954 104058 181986 104294
rect 182222 104058 182306 104294
rect 182542 104058 182574 104294
rect 181954 68614 182574 104058
rect 181954 68378 181986 68614
rect 182222 68378 182306 68614
rect 182542 68378 182574 68614
rect 181954 68294 182574 68378
rect 181954 68058 181986 68294
rect 182222 68058 182306 68294
rect 182542 68058 182574 68294
rect 181954 32614 182574 68058
rect 181954 32378 181986 32614
rect 182222 32378 182306 32614
rect 182542 32378 182574 32614
rect 181954 32294 182574 32378
rect 181954 32058 181986 32294
rect 182222 32058 182306 32294
rect 182542 32058 182574 32294
rect 178234 -5382 178266 -5146
rect 178502 -5382 178586 -5146
rect 178822 -5382 178854 -5146
rect 178234 -5466 178854 -5382
rect 178234 -5702 178266 -5466
rect 178502 -5702 178586 -5466
rect 178822 -5702 178854 -5466
rect 178234 -5734 178854 -5702
rect 171954 -6342 171986 -6106
rect 172222 -6342 172306 -6106
rect 172542 -6342 172574 -6106
rect 171954 -6426 172574 -6342
rect 171954 -6662 171986 -6426
rect 172222 -6662 172306 -6426
rect 172542 -6662 172574 -6426
rect 171954 -7654 172574 -6662
rect 181954 -7066 182574 32058
rect 184514 706758 185134 707750
rect 184514 706522 184546 706758
rect 184782 706522 184866 706758
rect 185102 706522 185134 706758
rect 184514 706438 185134 706522
rect 184514 706202 184546 706438
rect 184782 706202 184866 706438
rect 185102 706202 185134 706438
rect 184514 691174 185134 706202
rect 184514 690938 184546 691174
rect 184782 690938 184866 691174
rect 185102 690938 185134 691174
rect 184514 690854 185134 690938
rect 184514 690618 184546 690854
rect 184782 690618 184866 690854
rect 185102 690618 185134 690854
rect 184514 655174 185134 690618
rect 184514 654938 184546 655174
rect 184782 654938 184866 655174
rect 185102 654938 185134 655174
rect 184514 654854 185134 654938
rect 184514 654618 184546 654854
rect 184782 654618 184866 654854
rect 185102 654618 185134 654854
rect 184514 619174 185134 654618
rect 184514 618938 184546 619174
rect 184782 618938 184866 619174
rect 185102 618938 185134 619174
rect 184514 618854 185134 618938
rect 184514 618618 184546 618854
rect 184782 618618 184866 618854
rect 185102 618618 185134 618854
rect 184514 583174 185134 618618
rect 184514 582938 184546 583174
rect 184782 582938 184866 583174
rect 185102 582938 185134 583174
rect 184514 582854 185134 582938
rect 184514 582618 184546 582854
rect 184782 582618 184866 582854
rect 185102 582618 185134 582854
rect 184514 547174 185134 582618
rect 184514 546938 184546 547174
rect 184782 546938 184866 547174
rect 185102 546938 185134 547174
rect 184514 546854 185134 546938
rect 184514 546618 184546 546854
rect 184782 546618 184866 546854
rect 185102 546618 185134 546854
rect 184514 511174 185134 546618
rect 184514 510938 184546 511174
rect 184782 510938 184866 511174
rect 185102 510938 185134 511174
rect 184514 510854 185134 510938
rect 184514 510618 184546 510854
rect 184782 510618 184866 510854
rect 185102 510618 185134 510854
rect 184514 475174 185134 510618
rect 184514 474938 184546 475174
rect 184782 474938 184866 475174
rect 185102 474938 185134 475174
rect 184514 474854 185134 474938
rect 184514 474618 184546 474854
rect 184782 474618 184866 474854
rect 185102 474618 185134 474854
rect 184514 439174 185134 474618
rect 184514 438938 184546 439174
rect 184782 438938 184866 439174
rect 185102 438938 185134 439174
rect 184514 438854 185134 438938
rect 184514 438618 184546 438854
rect 184782 438618 184866 438854
rect 185102 438618 185134 438854
rect 184514 403174 185134 438618
rect 184514 402938 184546 403174
rect 184782 402938 184866 403174
rect 185102 402938 185134 403174
rect 184514 402854 185134 402938
rect 184514 402618 184546 402854
rect 184782 402618 184866 402854
rect 185102 402618 185134 402854
rect 184514 367174 185134 402618
rect 184514 366938 184546 367174
rect 184782 366938 184866 367174
rect 185102 366938 185134 367174
rect 184514 366854 185134 366938
rect 184514 366618 184546 366854
rect 184782 366618 184866 366854
rect 185102 366618 185134 366854
rect 184514 331174 185134 366618
rect 184514 330938 184546 331174
rect 184782 330938 184866 331174
rect 185102 330938 185134 331174
rect 184514 330854 185134 330938
rect 184514 330618 184546 330854
rect 184782 330618 184866 330854
rect 185102 330618 185134 330854
rect 184514 295174 185134 330618
rect 184514 294938 184546 295174
rect 184782 294938 184866 295174
rect 185102 294938 185134 295174
rect 184514 294854 185134 294938
rect 184514 294618 184546 294854
rect 184782 294618 184866 294854
rect 185102 294618 185134 294854
rect 184514 259174 185134 294618
rect 184514 258938 184546 259174
rect 184782 258938 184866 259174
rect 185102 258938 185134 259174
rect 184514 258854 185134 258938
rect 184514 258618 184546 258854
rect 184782 258618 184866 258854
rect 185102 258618 185134 258854
rect 184514 223174 185134 258618
rect 184514 222938 184546 223174
rect 184782 222938 184866 223174
rect 185102 222938 185134 223174
rect 184514 222854 185134 222938
rect 184514 222618 184546 222854
rect 184782 222618 184866 222854
rect 185102 222618 185134 222854
rect 184514 187174 185134 222618
rect 184514 186938 184546 187174
rect 184782 186938 184866 187174
rect 185102 186938 185134 187174
rect 184514 186854 185134 186938
rect 184514 186618 184546 186854
rect 184782 186618 184866 186854
rect 185102 186618 185134 186854
rect 184514 151174 185134 186618
rect 184514 150938 184546 151174
rect 184782 150938 184866 151174
rect 185102 150938 185134 151174
rect 184514 150854 185134 150938
rect 184514 150618 184546 150854
rect 184782 150618 184866 150854
rect 185102 150618 185134 150854
rect 184514 115174 185134 150618
rect 184514 114938 184546 115174
rect 184782 114938 184866 115174
rect 185102 114938 185134 115174
rect 184514 114854 185134 114938
rect 184514 114618 184546 114854
rect 184782 114618 184866 114854
rect 185102 114618 185134 114854
rect 184514 79174 185134 114618
rect 184514 78938 184546 79174
rect 184782 78938 184866 79174
rect 185102 78938 185134 79174
rect 184514 78854 185134 78938
rect 184514 78618 184546 78854
rect 184782 78618 184866 78854
rect 185102 78618 185134 78854
rect 184514 43174 185134 78618
rect 184514 42938 184546 43174
rect 184782 42938 184866 43174
rect 185102 42938 185134 43174
rect 184514 42854 185134 42938
rect 184514 42618 184546 42854
rect 184782 42618 184866 42854
rect 185102 42618 185134 42854
rect 184514 7174 185134 42618
rect 184514 6938 184546 7174
rect 184782 6938 184866 7174
rect 185102 6938 185134 7174
rect 184514 6854 185134 6938
rect 184514 6618 184546 6854
rect 184782 6618 184866 6854
rect 185102 6618 185134 6854
rect 184514 -2266 185134 6618
rect 184514 -2502 184546 -2266
rect 184782 -2502 184866 -2266
rect 185102 -2502 185134 -2266
rect 184514 -2586 185134 -2502
rect 184514 -2822 184546 -2586
rect 184782 -2822 184866 -2586
rect 185102 -2822 185134 -2586
rect 184514 -3814 185134 -2822
rect 188234 694894 188854 708122
rect 188234 694658 188266 694894
rect 188502 694658 188586 694894
rect 188822 694658 188854 694894
rect 188234 694574 188854 694658
rect 188234 694338 188266 694574
rect 188502 694338 188586 694574
rect 188822 694338 188854 694574
rect 188234 658894 188854 694338
rect 188234 658658 188266 658894
rect 188502 658658 188586 658894
rect 188822 658658 188854 658894
rect 188234 658574 188854 658658
rect 188234 658338 188266 658574
rect 188502 658338 188586 658574
rect 188822 658338 188854 658574
rect 188234 622894 188854 658338
rect 188234 622658 188266 622894
rect 188502 622658 188586 622894
rect 188822 622658 188854 622894
rect 188234 622574 188854 622658
rect 188234 622338 188266 622574
rect 188502 622338 188586 622574
rect 188822 622338 188854 622574
rect 188234 586894 188854 622338
rect 188234 586658 188266 586894
rect 188502 586658 188586 586894
rect 188822 586658 188854 586894
rect 188234 586574 188854 586658
rect 188234 586338 188266 586574
rect 188502 586338 188586 586574
rect 188822 586338 188854 586574
rect 188234 550894 188854 586338
rect 188234 550658 188266 550894
rect 188502 550658 188586 550894
rect 188822 550658 188854 550894
rect 188234 550574 188854 550658
rect 188234 550338 188266 550574
rect 188502 550338 188586 550574
rect 188822 550338 188854 550574
rect 188234 514894 188854 550338
rect 188234 514658 188266 514894
rect 188502 514658 188586 514894
rect 188822 514658 188854 514894
rect 188234 514574 188854 514658
rect 188234 514338 188266 514574
rect 188502 514338 188586 514574
rect 188822 514338 188854 514574
rect 188234 478894 188854 514338
rect 188234 478658 188266 478894
rect 188502 478658 188586 478894
rect 188822 478658 188854 478894
rect 188234 478574 188854 478658
rect 188234 478338 188266 478574
rect 188502 478338 188586 478574
rect 188822 478338 188854 478574
rect 188234 442894 188854 478338
rect 188234 442658 188266 442894
rect 188502 442658 188586 442894
rect 188822 442658 188854 442894
rect 188234 442574 188854 442658
rect 188234 442338 188266 442574
rect 188502 442338 188586 442574
rect 188822 442338 188854 442574
rect 188234 406894 188854 442338
rect 188234 406658 188266 406894
rect 188502 406658 188586 406894
rect 188822 406658 188854 406894
rect 188234 406574 188854 406658
rect 188234 406338 188266 406574
rect 188502 406338 188586 406574
rect 188822 406338 188854 406574
rect 188234 370894 188854 406338
rect 188234 370658 188266 370894
rect 188502 370658 188586 370894
rect 188822 370658 188854 370894
rect 188234 370574 188854 370658
rect 188234 370338 188266 370574
rect 188502 370338 188586 370574
rect 188822 370338 188854 370574
rect 188234 334894 188854 370338
rect 188234 334658 188266 334894
rect 188502 334658 188586 334894
rect 188822 334658 188854 334894
rect 188234 334574 188854 334658
rect 188234 334338 188266 334574
rect 188502 334338 188586 334574
rect 188822 334338 188854 334574
rect 188234 298894 188854 334338
rect 188234 298658 188266 298894
rect 188502 298658 188586 298894
rect 188822 298658 188854 298894
rect 188234 298574 188854 298658
rect 188234 298338 188266 298574
rect 188502 298338 188586 298574
rect 188822 298338 188854 298574
rect 188234 262894 188854 298338
rect 188234 262658 188266 262894
rect 188502 262658 188586 262894
rect 188822 262658 188854 262894
rect 188234 262574 188854 262658
rect 188234 262338 188266 262574
rect 188502 262338 188586 262574
rect 188822 262338 188854 262574
rect 188234 226894 188854 262338
rect 188234 226658 188266 226894
rect 188502 226658 188586 226894
rect 188822 226658 188854 226894
rect 188234 226574 188854 226658
rect 188234 226338 188266 226574
rect 188502 226338 188586 226574
rect 188822 226338 188854 226574
rect 188234 190894 188854 226338
rect 188234 190658 188266 190894
rect 188502 190658 188586 190894
rect 188822 190658 188854 190894
rect 188234 190574 188854 190658
rect 188234 190338 188266 190574
rect 188502 190338 188586 190574
rect 188822 190338 188854 190574
rect 188234 154894 188854 190338
rect 188234 154658 188266 154894
rect 188502 154658 188586 154894
rect 188822 154658 188854 154894
rect 188234 154574 188854 154658
rect 188234 154338 188266 154574
rect 188502 154338 188586 154574
rect 188822 154338 188854 154574
rect 188234 118894 188854 154338
rect 188234 118658 188266 118894
rect 188502 118658 188586 118894
rect 188822 118658 188854 118894
rect 188234 118574 188854 118658
rect 188234 118338 188266 118574
rect 188502 118338 188586 118574
rect 188822 118338 188854 118574
rect 188234 82894 188854 118338
rect 188234 82658 188266 82894
rect 188502 82658 188586 82894
rect 188822 82658 188854 82894
rect 188234 82574 188854 82658
rect 188234 82338 188266 82574
rect 188502 82338 188586 82574
rect 188822 82338 188854 82574
rect 188234 46894 188854 82338
rect 188234 46658 188266 46894
rect 188502 46658 188586 46894
rect 188822 46658 188854 46894
rect 188234 46574 188854 46658
rect 188234 46338 188266 46574
rect 188502 46338 188586 46574
rect 188822 46338 188854 46574
rect 188234 10894 188854 46338
rect 188234 10658 188266 10894
rect 188502 10658 188586 10894
rect 188822 10658 188854 10894
rect 188234 10574 188854 10658
rect 188234 10338 188266 10574
rect 188502 10338 188586 10574
rect 188822 10338 188854 10574
rect 188234 -4186 188854 10338
rect 190794 705798 191414 705830
rect 190794 705562 190826 705798
rect 191062 705562 191146 705798
rect 191382 705562 191414 705798
rect 190794 705478 191414 705562
rect 190794 705242 190826 705478
rect 191062 705242 191146 705478
rect 191382 705242 191414 705478
rect 190794 669454 191414 705242
rect 190794 669218 190826 669454
rect 191062 669218 191146 669454
rect 191382 669218 191414 669454
rect 190794 669134 191414 669218
rect 190794 668898 190826 669134
rect 191062 668898 191146 669134
rect 191382 668898 191414 669134
rect 190794 633454 191414 668898
rect 190794 633218 190826 633454
rect 191062 633218 191146 633454
rect 191382 633218 191414 633454
rect 190794 633134 191414 633218
rect 190794 632898 190826 633134
rect 191062 632898 191146 633134
rect 191382 632898 191414 633134
rect 190794 597454 191414 632898
rect 190794 597218 190826 597454
rect 191062 597218 191146 597454
rect 191382 597218 191414 597454
rect 190794 597134 191414 597218
rect 190794 596898 190826 597134
rect 191062 596898 191146 597134
rect 191382 596898 191414 597134
rect 190794 561454 191414 596898
rect 190794 561218 190826 561454
rect 191062 561218 191146 561454
rect 191382 561218 191414 561454
rect 190794 561134 191414 561218
rect 190794 560898 190826 561134
rect 191062 560898 191146 561134
rect 191382 560898 191414 561134
rect 190794 525454 191414 560898
rect 190794 525218 190826 525454
rect 191062 525218 191146 525454
rect 191382 525218 191414 525454
rect 190794 525134 191414 525218
rect 190794 524898 190826 525134
rect 191062 524898 191146 525134
rect 191382 524898 191414 525134
rect 190794 489454 191414 524898
rect 190794 489218 190826 489454
rect 191062 489218 191146 489454
rect 191382 489218 191414 489454
rect 190794 489134 191414 489218
rect 190794 488898 190826 489134
rect 191062 488898 191146 489134
rect 191382 488898 191414 489134
rect 190794 453454 191414 488898
rect 190794 453218 190826 453454
rect 191062 453218 191146 453454
rect 191382 453218 191414 453454
rect 190794 453134 191414 453218
rect 190794 452898 190826 453134
rect 191062 452898 191146 453134
rect 191382 452898 191414 453134
rect 190794 417454 191414 452898
rect 190794 417218 190826 417454
rect 191062 417218 191146 417454
rect 191382 417218 191414 417454
rect 190794 417134 191414 417218
rect 190794 416898 190826 417134
rect 191062 416898 191146 417134
rect 191382 416898 191414 417134
rect 190794 381454 191414 416898
rect 190794 381218 190826 381454
rect 191062 381218 191146 381454
rect 191382 381218 191414 381454
rect 190794 381134 191414 381218
rect 190794 380898 190826 381134
rect 191062 380898 191146 381134
rect 191382 380898 191414 381134
rect 190794 345454 191414 380898
rect 190794 345218 190826 345454
rect 191062 345218 191146 345454
rect 191382 345218 191414 345454
rect 190794 345134 191414 345218
rect 190794 344898 190826 345134
rect 191062 344898 191146 345134
rect 191382 344898 191414 345134
rect 190794 309454 191414 344898
rect 190794 309218 190826 309454
rect 191062 309218 191146 309454
rect 191382 309218 191414 309454
rect 190794 309134 191414 309218
rect 190794 308898 190826 309134
rect 191062 308898 191146 309134
rect 191382 308898 191414 309134
rect 190794 273454 191414 308898
rect 190794 273218 190826 273454
rect 191062 273218 191146 273454
rect 191382 273218 191414 273454
rect 190794 273134 191414 273218
rect 190794 272898 190826 273134
rect 191062 272898 191146 273134
rect 191382 272898 191414 273134
rect 190794 237454 191414 272898
rect 190794 237218 190826 237454
rect 191062 237218 191146 237454
rect 191382 237218 191414 237454
rect 190794 237134 191414 237218
rect 190794 236898 190826 237134
rect 191062 236898 191146 237134
rect 191382 236898 191414 237134
rect 190794 201454 191414 236898
rect 190794 201218 190826 201454
rect 191062 201218 191146 201454
rect 191382 201218 191414 201454
rect 190794 201134 191414 201218
rect 190794 200898 190826 201134
rect 191062 200898 191146 201134
rect 191382 200898 191414 201134
rect 190794 165454 191414 200898
rect 190794 165218 190826 165454
rect 191062 165218 191146 165454
rect 191382 165218 191414 165454
rect 190794 165134 191414 165218
rect 190794 164898 190826 165134
rect 191062 164898 191146 165134
rect 191382 164898 191414 165134
rect 190794 129454 191414 164898
rect 190794 129218 190826 129454
rect 191062 129218 191146 129454
rect 191382 129218 191414 129454
rect 190794 129134 191414 129218
rect 190794 128898 190826 129134
rect 191062 128898 191146 129134
rect 191382 128898 191414 129134
rect 190794 93454 191414 128898
rect 190794 93218 190826 93454
rect 191062 93218 191146 93454
rect 191382 93218 191414 93454
rect 190794 93134 191414 93218
rect 190794 92898 190826 93134
rect 191062 92898 191146 93134
rect 191382 92898 191414 93134
rect 190794 57454 191414 92898
rect 190794 57218 190826 57454
rect 191062 57218 191146 57454
rect 191382 57218 191414 57454
rect 190794 57134 191414 57218
rect 190794 56898 190826 57134
rect 191062 56898 191146 57134
rect 191382 56898 191414 57134
rect 190794 21454 191414 56898
rect 190794 21218 190826 21454
rect 191062 21218 191146 21454
rect 191382 21218 191414 21454
rect 190794 21134 191414 21218
rect 190794 20898 190826 21134
rect 191062 20898 191146 21134
rect 191382 20898 191414 21134
rect 190794 -1306 191414 20898
rect 190794 -1542 190826 -1306
rect 191062 -1542 191146 -1306
rect 191382 -1542 191414 -1306
rect 190794 -1626 191414 -1542
rect 190794 -1862 190826 -1626
rect 191062 -1862 191146 -1626
rect 191382 -1862 191414 -1626
rect 190794 -1894 191414 -1862
rect 191954 698614 192574 710042
rect 201954 711558 202574 711590
rect 201954 711322 201986 711558
rect 202222 711322 202306 711558
rect 202542 711322 202574 711558
rect 201954 711238 202574 711322
rect 201954 711002 201986 711238
rect 202222 711002 202306 711238
rect 202542 711002 202574 711238
rect 198234 709638 198854 709670
rect 198234 709402 198266 709638
rect 198502 709402 198586 709638
rect 198822 709402 198854 709638
rect 198234 709318 198854 709402
rect 198234 709082 198266 709318
rect 198502 709082 198586 709318
rect 198822 709082 198854 709318
rect 191954 698378 191986 698614
rect 192222 698378 192306 698614
rect 192542 698378 192574 698614
rect 191954 698294 192574 698378
rect 191954 698058 191986 698294
rect 192222 698058 192306 698294
rect 192542 698058 192574 698294
rect 191954 662614 192574 698058
rect 191954 662378 191986 662614
rect 192222 662378 192306 662614
rect 192542 662378 192574 662614
rect 191954 662294 192574 662378
rect 191954 662058 191986 662294
rect 192222 662058 192306 662294
rect 192542 662058 192574 662294
rect 191954 626614 192574 662058
rect 191954 626378 191986 626614
rect 192222 626378 192306 626614
rect 192542 626378 192574 626614
rect 191954 626294 192574 626378
rect 191954 626058 191986 626294
rect 192222 626058 192306 626294
rect 192542 626058 192574 626294
rect 191954 590614 192574 626058
rect 191954 590378 191986 590614
rect 192222 590378 192306 590614
rect 192542 590378 192574 590614
rect 191954 590294 192574 590378
rect 191954 590058 191986 590294
rect 192222 590058 192306 590294
rect 192542 590058 192574 590294
rect 191954 554614 192574 590058
rect 191954 554378 191986 554614
rect 192222 554378 192306 554614
rect 192542 554378 192574 554614
rect 191954 554294 192574 554378
rect 191954 554058 191986 554294
rect 192222 554058 192306 554294
rect 192542 554058 192574 554294
rect 191954 518614 192574 554058
rect 191954 518378 191986 518614
rect 192222 518378 192306 518614
rect 192542 518378 192574 518614
rect 191954 518294 192574 518378
rect 191954 518058 191986 518294
rect 192222 518058 192306 518294
rect 192542 518058 192574 518294
rect 191954 482614 192574 518058
rect 191954 482378 191986 482614
rect 192222 482378 192306 482614
rect 192542 482378 192574 482614
rect 191954 482294 192574 482378
rect 191954 482058 191986 482294
rect 192222 482058 192306 482294
rect 192542 482058 192574 482294
rect 191954 446614 192574 482058
rect 191954 446378 191986 446614
rect 192222 446378 192306 446614
rect 192542 446378 192574 446614
rect 191954 446294 192574 446378
rect 191954 446058 191986 446294
rect 192222 446058 192306 446294
rect 192542 446058 192574 446294
rect 191954 410614 192574 446058
rect 191954 410378 191986 410614
rect 192222 410378 192306 410614
rect 192542 410378 192574 410614
rect 191954 410294 192574 410378
rect 191954 410058 191986 410294
rect 192222 410058 192306 410294
rect 192542 410058 192574 410294
rect 191954 374614 192574 410058
rect 191954 374378 191986 374614
rect 192222 374378 192306 374614
rect 192542 374378 192574 374614
rect 191954 374294 192574 374378
rect 191954 374058 191986 374294
rect 192222 374058 192306 374294
rect 192542 374058 192574 374294
rect 191954 338614 192574 374058
rect 191954 338378 191986 338614
rect 192222 338378 192306 338614
rect 192542 338378 192574 338614
rect 191954 338294 192574 338378
rect 191954 338058 191986 338294
rect 192222 338058 192306 338294
rect 192542 338058 192574 338294
rect 191954 302614 192574 338058
rect 191954 302378 191986 302614
rect 192222 302378 192306 302614
rect 192542 302378 192574 302614
rect 191954 302294 192574 302378
rect 191954 302058 191986 302294
rect 192222 302058 192306 302294
rect 192542 302058 192574 302294
rect 191954 266614 192574 302058
rect 191954 266378 191986 266614
rect 192222 266378 192306 266614
rect 192542 266378 192574 266614
rect 191954 266294 192574 266378
rect 191954 266058 191986 266294
rect 192222 266058 192306 266294
rect 192542 266058 192574 266294
rect 191954 230614 192574 266058
rect 191954 230378 191986 230614
rect 192222 230378 192306 230614
rect 192542 230378 192574 230614
rect 191954 230294 192574 230378
rect 191954 230058 191986 230294
rect 192222 230058 192306 230294
rect 192542 230058 192574 230294
rect 191954 194614 192574 230058
rect 191954 194378 191986 194614
rect 192222 194378 192306 194614
rect 192542 194378 192574 194614
rect 191954 194294 192574 194378
rect 191954 194058 191986 194294
rect 192222 194058 192306 194294
rect 192542 194058 192574 194294
rect 191954 158614 192574 194058
rect 191954 158378 191986 158614
rect 192222 158378 192306 158614
rect 192542 158378 192574 158614
rect 191954 158294 192574 158378
rect 191954 158058 191986 158294
rect 192222 158058 192306 158294
rect 192542 158058 192574 158294
rect 191954 122614 192574 158058
rect 191954 122378 191986 122614
rect 192222 122378 192306 122614
rect 192542 122378 192574 122614
rect 191954 122294 192574 122378
rect 191954 122058 191986 122294
rect 192222 122058 192306 122294
rect 192542 122058 192574 122294
rect 191954 86614 192574 122058
rect 191954 86378 191986 86614
rect 192222 86378 192306 86614
rect 192542 86378 192574 86614
rect 191954 86294 192574 86378
rect 191954 86058 191986 86294
rect 192222 86058 192306 86294
rect 192542 86058 192574 86294
rect 191954 50614 192574 86058
rect 191954 50378 191986 50614
rect 192222 50378 192306 50614
rect 192542 50378 192574 50614
rect 191954 50294 192574 50378
rect 191954 50058 191986 50294
rect 192222 50058 192306 50294
rect 192542 50058 192574 50294
rect 191954 14614 192574 50058
rect 191954 14378 191986 14614
rect 192222 14378 192306 14614
rect 192542 14378 192574 14614
rect 191954 14294 192574 14378
rect 191954 14058 191986 14294
rect 192222 14058 192306 14294
rect 192542 14058 192574 14294
rect 188234 -4422 188266 -4186
rect 188502 -4422 188586 -4186
rect 188822 -4422 188854 -4186
rect 188234 -4506 188854 -4422
rect 188234 -4742 188266 -4506
rect 188502 -4742 188586 -4506
rect 188822 -4742 188854 -4506
rect 188234 -5734 188854 -4742
rect 181954 -7302 181986 -7066
rect 182222 -7302 182306 -7066
rect 182542 -7302 182574 -7066
rect 181954 -7386 182574 -7302
rect 181954 -7622 181986 -7386
rect 182222 -7622 182306 -7386
rect 182542 -7622 182574 -7386
rect 181954 -7654 182574 -7622
rect 191954 -6106 192574 14058
rect 194514 707718 195134 707750
rect 194514 707482 194546 707718
rect 194782 707482 194866 707718
rect 195102 707482 195134 707718
rect 194514 707398 195134 707482
rect 194514 707162 194546 707398
rect 194782 707162 194866 707398
rect 195102 707162 195134 707398
rect 194514 673174 195134 707162
rect 194514 672938 194546 673174
rect 194782 672938 194866 673174
rect 195102 672938 195134 673174
rect 194514 672854 195134 672938
rect 194514 672618 194546 672854
rect 194782 672618 194866 672854
rect 195102 672618 195134 672854
rect 194514 637174 195134 672618
rect 194514 636938 194546 637174
rect 194782 636938 194866 637174
rect 195102 636938 195134 637174
rect 194514 636854 195134 636938
rect 194514 636618 194546 636854
rect 194782 636618 194866 636854
rect 195102 636618 195134 636854
rect 194514 601174 195134 636618
rect 194514 600938 194546 601174
rect 194782 600938 194866 601174
rect 195102 600938 195134 601174
rect 194514 600854 195134 600938
rect 194514 600618 194546 600854
rect 194782 600618 194866 600854
rect 195102 600618 195134 600854
rect 194514 565174 195134 600618
rect 194514 564938 194546 565174
rect 194782 564938 194866 565174
rect 195102 564938 195134 565174
rect 194514 564854 195134 564938
rect 194514 564618 194546 564854
rect 194782 564618 194866 564854
rect 195102 564618 195134 564854
rect 194514 529174 195134 564618
rect 194514 528938 194546 529174
rect 194782 528938 194866 529174
rect 195102 528938 195134 529174
rect 194514 528854 195134 528938
rect 194514 528618 194546 528854
rect 194782 528618 194866 528854
rect 195102 528618 195134 528854
rect 194514 493174 195134 528618
rect 194514 492938 194546 493174
rect 194782 492938 194866 493174
rect 195102 492938 195134 493174
rect 194514 492854 195134 492938
rect 194514 492618 194546 492854
rect 194782 492618 194866 492854
rect 195102 492618 195134 492854
rect 194514 457174 195134 492618
rect 194514 456938 194546 457174
rect 194782 456938 194866 457174
rect 195102 456938 195134 457174
rect 194514 456854 195134 456938
rect 194514 456618 194546 456854
rect 194782 456618 194866 456854
rect 195102 456618 195134 456854
rect 194514 421174 195134 456618
rect 194514 420938 194546 421174
rect 194782 420938 194866 421174
rect 195102 420938 195134 421174
rect 194514 420854 195134 420938
rect 194514 420618 194546 420854
rect 194782 420618 194866 420854
rect 195102 420618 195134 420854
rect 194514 385174 195134 420618
rect 194514 384938 194546 385174
rect 194782 384938 194866 385174
rect 195102 384938 195134 385174
rect 194514 384854 195134 384938
rect 194514 384618 194546 384854
rect 194782 384618 194866 384854
rect 195102 384618 195134 384854
rect 194514 349174 195134 384618
rect 194514 348938 194546 349174
rect 194782 348938 194866 349174
rect 195102 348938 195134 349174
rect 194514 348854 195134 348938
rect 194514 348618 194546 348854
rect 194782 348618 194866 348854
rect 195102 348618 195134 348854
rect 194514 313174 195134 348618
rect 194514 312938 194546 313174
rect 194782 312938 194866 313174
rect 195102 312938 195134 313174
rect 194514 312854 195134 312938
rect 194514 312618 194546 312854
rect 194782 312618 194866 312854
rect 195102 312618 195134 312854
rect 194514 277174 195134 312618
rect 194514 276938 194546 277174
rect 194782 276938 194866 277174
rect 195102 276938 195134 277174
rect 194514 276854 195134 276938
rect 194514 276618 194546 276854
rect 194782 276618 194866 276854
rect 195102 276618 195134 276854
rect 194514 241174 195134 276618
rect 194514 240938 194546 241174
rect 194782 240938 194866 241174
rect 195102 240938 195134 241174
rect 194514 240854 195134 240938
rect 194514 240618 194546 240854
rect 194782 240618 194866 240854
rect 195102 240618 195134 240854
rect 194514 205174 195134 240618
rect 194514 204938 194546 205174
rect 194782 204938 194866 205174
rect 195102 204938 195134 205174
rect 194514 204854 195134 204938
rect 194514 204618 194546 204854
rect 194782 204618 194866 204854
rect 195102 204618 195134 204854
rect 194514 169174 195134 204618
rect 194514 168938 194546 169174
rect 194782 168938 194866 169174
rect 195102 168938 195134 169174
rect 194514 168854 195134 168938
rect 194514 168618 194546 168854
rect 194782 168618 194866 168854
rect 195102 168618 195134 168854
rect 194514 133174 195134 168618
rect 194514 132938 194546 133174
rect 194782 132938 194866 133174
rect 195102 132938 195134 133174
rect 194514 132854 195134 132938
rect 194514 132618 194546 132854
rect 194782 132618 194866 132854
rect 195102 132618 195134 132854
rect 194514 97174 195134 132618
rect 194514 96938 194546 97174
rect 194782 96938 194866 97174
rect 195102 96938 195134 97174
rect 194514 96854 195134 96938
rect 194514 96618 194546 96854
rect 194782 96618 194866 96854
rect 195102 96618 195134 96854
rect 194514 61174 195134 96618
rect 194514 60938 194546 61174
rect 194782 60938 194866 61174
rect 195102 60938 195134 61174
rect 194514 60854 195134 60938
rect 194514 60618 194546 60854
rect 194782 60618 194866 60854
rect 195102 60618 195134 60854
rect 194514 25174 195134 60618
rect 194514 24938 194546 25174
rect 194782 24938 194866 25174
rect 195102 24938 195134 25174
rect 194514 24854 195134 24938
rect 194514 24618 194546 24854
rect 194782 24618 194866 24854
rect 195102 24618 195134 24854
rect 194514 -3226 195134 24618
rect 194514 -3462 194546 -3226
rect 194782 -3462 194866 -3226
rect 195102 -3462 195134 -3226
rect 194514 -3546 195134 -3462
rect 194514 -3782 194546 -3546
rect 194782 -3782 194866 -3546
rect 195102 -3782 195134 -3546
rect 194514 -3814 195134 -3782
rect 198234 676894 198854 709082
rect 198234 676658 198266 676894
rect 198502 676658 198586 676894
rect 198822 676658 198854 676894
rect 198234 676574 198854 676658
rect 198234 676338 198266 676574
rect 198502 676338 198586 676574
rect 198822 676338 198854 676574
rect 198234 640894 198854 676338
rect 198234 640658 198266 640894
rect 198502 640658 198586 640894
rect 198822 640658 198854 640894
rect 198234 640574 198854 640658
rect 198234 640338 198266 640574
rect 198502 640338 198586 640574
rect 198822 640338 198854 640574
rect 198234 604894 198854 640338
rect 198234 604658 198266 604894
rect 198502 604658 198586 604894
rect 198822 604658 198854 604894
rect 198234 604574 198854 604658
rect 198234 604338 198266 604574
rect 198502 604338 198586 604574
rect 198822 604338 198854 604574
rect 198234 568894 198854 604338
rect 198234 568658 198266 568894
rect 198502 568658 198586 568894
rect 198822 568658 198854 568894
rect 198234 568574 198854 568658
rect 198234 568338 198266 568574
rect 198502 568338 198586 568574
rect 198822 568338 198854 568574
rect 198234 532894 198854 568338
rect 198234 532658 198266 532894
rect 198502 532658 198586 532894
rect 198822 532658 198854 532894
rect 198234 532574 198854 532658
rect 198234 532338 198266 532574
rect 198502 532338 198586 532574
rect 198822 532338 198854 532574
rect 198234 496894 198854 532338
rect 198234 496658 198266 496894
rect 198502 496658 198586 496894
rect 198822 496658 198854 496894
rect 198234 496574 198854 496658
rect 198234 496338 198266 496574
rect 198502 496338 198586 496574
rect 198822 496338 198854 496574
rect 198234 460894 198854 496338
rect 198234 460658 198266 460894
rect 198502 460658 198586 460894
rect 198822 460658 198854 460894
rect 198234 460574 198854 460658
rect 198234 460338 198266 460574
rect 198502 460338 198586 460574
rect 198822 460338 198854 460574
rect 198234 424894 198854 460338
rect 198234 424658 198266 424894
rect 198502 424658 198586 424894
rect 198822 424658 198854 424894
rect 198234 424574 198854 424658
rect 198234 424338 198266 424574
rect 198502 424338 198586 424574
rect 198822 424338 198854 424574
rect 198234 388894 198854 424338
rect 198234 388658 198266 388894
rect 198502 388658 198586 388894
rect 198822 388658 198854 388894
rect 198234 388574 198854 388658
rect 198234 388338 198266 388574
rect 198502 388338 198586 388574
rect 198822 388338 198854 388574
rect 198234 352894 198854 388338
rect 198234 352658 198266 352894
rect 198502 352658 198586 352894
rect 198822 352658 198854 352894
rect 198234 352574 198854 352658
rect 198234 352338 198266 352574
rect 198502 352338 198586 352574
rect 198822 352338 198854 352574
rect 198234 316894 198854 352338
rect 198234 316658 198266 316894
rect 198502 316658 198586 316894
rect 198822 316658 198854 316894
rect 198234 316574 198854 316658
rect 198234 316338 198266 316574
rect 198502 316338 198586 316574
rect 198822 316338 198854 316574
rect 198234 280894 198854 316338
rect 198234 280658 198266 280894
rect 198502 280658 198586 280894
rect 198822 280658 198854 280894
rect 198234 280574 198854 280658
rect 198234 280338 198266 280574
rect 198502 280338 198586 280574
rect 198822 280338 198854 280574
rect 198234 244894 198854 280338
rect 198234 244658 198266 244894
rect 198502 244658 198586 244894
rect 198822 244658 198854 244894
rect 198234 244574 198854 244658
rect 198234 244338 198266 244574
rect 198502 244338 198586 244574
rect 198822 244338 198854 244574
rect 198234 208894 198854 244338
rect 198234 208658 198266 208894
rect 198502 208658 198586 208894
rect 198822 208658 198854 208894
rect 198234 208574 198854 208658
rect 198234 208338 198266 208574
rect 198502 208338 198586 208574
rect 198822 208338 198854 208574
rect 198234 172894 198854 208338
rect 198234 172658 198266 172894
rect 198502 172658 198586 172894
rect 198822 172658 198854 172894
rect 198234 172574 198854 172658
rect 198234 172338 198266 172574
rect 198502 172338 198586 172574
rect 198822 172338 198854 172574
rect 198234 136894 198854 172338
rect 198234 136658 198266 136894
rect 198502 136658 198586 136894
rect 198822 136658 198854 136894
rect 198234 136574 198854 136658
rect 198234 136338 198266 136574
rect 198502 136338 198586 136574
rect 198822 136338 198854 136574
rect 198234 100894 198854 136338
rect 198234 100658 198266 100894
rect 198502 100658 198586 100894
rect 198822 100658 198854 100894
rect 198234 100574 198854 100658
rect 198234 100338 198266 100574
rect 198502 100338 198586 100574
rect 198822 100338 198854 100574
rect 198234 64894 198854 100338
rect 198234 64658 198266 64894
rect 198502 64658 198586 64894
rect 198822 64658 198854 64894
rect 198234 64574 198854 64658
rect 198234 64338 198266 64574
rect 198502 64338 198586 64574
rect 198822 64338 198854 64574
rect 198234 28894 198854 64338
rect 198234 28658 198266 28894
rect 198502 28658 198586 28894
rect 198822 28658 198854 28894
rect 198234 28574 198854 28658
rect 198234 28338 198266 28574
rect 198502 28338 198586 28574
rect 198822 28338 198854 28574
rect 198234 -5146 198854 28338
rect 200794 704838 201414 705830
rect 200794 704602 200826 704838
rect 201062 704602 201146 704838
rect 201382 704602 201414 704838
rect 200794 704518 201414 704602
rect 200794 704282 200826 704518
rect 201062 704282 201146 704518
rect 201382 704282 201414 704518
rect 200794 687454 201414 704282
rect 200794 687218 200826 687454
rect 201062 687218 201146 687454
rect 201382 687218 201414 687454
rect 200794 687134 201414 687218
rect 200794 686898 200826 687134
rect 201062 686898 201146 687134
rect 201382 686898 201414 687134
rect 200794 651454 201414 686898
rect 200794 651218 200826 651454
rect 201062 651218 201146 651454
rect 201382 651218 201414 651454
rect 200794 651134 201414 651218
rect 200794 650898 200826 651134
rect 201062 650898 201146 651134
rect 201382 650898 201414 651134
rect 200794 615454 201414 650898
rect 200794 615218 200826 615454
rect 201062 615218 201146 615454
rect 201382 615218 201414 615454
rect 200794 615134 201414 615218
rect 200794 614898 200826 615134
rect 201062 614898 201146 615134
rect 201382 614898 201414 615134
rect 200794 579454 201414 614898
rect 200794 579218 200826 579454
rect 201062 579218 201146 579454
rect 201382 579218 201414 579454
rect 200794 579134 201414 579218
rect 200794 578898 200826 579134
rect 201062 578898 201146 579134
rect 201382 578898 201414 579134
rect 200794 543454 201414 578898
rect 200794 543218 200826 543454
rect 201062 543218 201146 543454
rect 201382 543218 201414 543454
rect 200794 543134 201414 543218
rect 200794 542898 200826 543134
rect 201062 542898 201146 543134
rect 201382 542898 201414 543134
rect 200794 507454 201414 542898
rect 200794 507218 200826 507454
rect 201062 507218 201146 507454
rect 201382 507218 201414 507454
rect 200794 507134 201414 507218
rect 200794 506898 200826 507134
rect 201062 506898 201146 507134
rect 201382 506898 201414 507134
rect 200794 471454 201414 506898
rect 200794 471218 200826 471454
rect 201062 471218 201146 471454
rect 201382 471218 201414 471454
rect 200794 471134 201414 471218
rect 200794 470898 200826 471134
rect 201062 470898 201146 471134
rect 201382 470898 201414 471134
rect 200794 435454 201414 470898
rect 200794 435218 200826 435454
rect 201062 435218 201146 435454
rect 201382 435218 201414 435454
rect 200794 435134 201414 435218
rect 200794 434898 200826 435134
rect 201062 434898 201146 435134
rect 201382 434898 201414 435134
rect 200794 399454 201414 434898
rect 200794 399218 200826 399454
rect 201062 399218 201146 399454
rect 201382 399218 201414 399454
rect 200794 399134 201414 399218
rect 200794 398898 200826 399134
rect 201062 398898 201146 399134
rect 201382 398898 201414 399134
rect 200794 363454 201414 398898
rect 200794 363218 200826 363454
rect 201062 363218 201146 363454
rect 201382 363218 201414 363454
rect 200794 363134 201414 363218
rect 200794 362898 200826 363134
rect 201062 362898 201146 363134
rect 201382 362898 201414 363134
rect 200794 327454 201414 362898
rect 200794 327218 200826 327454
rect 201062 327218 201146 327454
rect 201382 327218 201414 327454
rect 200794 327134 201414 327218
rect 200794 326898 200826 327134
rect 201062 326898 201146 327134
rect 201382 326898 201414 327134
rect 200794 291454 201414 326898
rect 200794 291218 200826 291454
rect 201062 291218 201146 291454
rect 201382 291218 201414 291454
rect 200794 291134 201414 291218
rect 200794 290898 200826 291134
rect 201062 290898 201146 291134
rect 201382 290898 201414 291134
rect 200794 255454 201414 290898
rect 200794 255218 200826 255454
rect 201062 255218 201146 255454
rect 201382 255218 201414 255454
rect 200794 255134 201414 255218
rect 200794 254898 200826 255134
rect 201062 254898 201146 255134
rect 201382 254898 201414 255134
rect 200794 219454 201414 254898
rect 200794 219218 200826 219454
rect 201062 219218 201146 219454
rect 201382 219218 201414 219454
rect 200794 219134 201414 219218
rect 200794 218898 200826 219134
rect 201062 218898 201146 219134
rect 201382 218898 201414 219134
rect 200794 183454 201414 218898
rect 200794 183218 200826 183454
rect 201062 183218 201146 183454
rect 201382 183218 201414 183454
rect 200794 183134 201414 183218
rect 200794 182898 200826 183134
rect 201062 182898 201146 183134
rect 201382 182898 201414 183134
rect 200794 147454 201414 182898
rect 200794 147218 200826 147454
rect 201062 147218 201146 147454
rect 201382 147218 201414 147454
rect 200794 147134 201414 147218
rect 200794 146898 200826 147134
rect 201062 146898 201146 147134
rect 201382 146898 201414 147134
rect 200794 111454 201414 146898
rect 200794 111218 200826 111454
rect 201062 111218 201146 111454
rect 201382 111218 201414 111454
rect 200794 111134 201414 111218
rect 200794 110898 200826 111134
rect 201062 110898 201146 111134
rect 201382 110898 201414 111134
rect 200794 75454 201414 110898
rect 200794 75218 200826 75454
rect 201062 75218 201146 75454
rect 201382 75218 201414 75454
rect 200794 75134 201414 75218
rect 200794 74898 200826 75134
rect 201062 74898 201146 75134
rect 201382 74898 201414 75134
rect 200794 39454 201414 74898
rect 200794 39218 200826 39454
rect 201062 39218 201146 39454
rect 201382 39218 201414 39454
rect 200794 39134 201414 39218
rect 200794 38898 200826 39134
rect 201062 38898 201146 39134
rect 201382 38898 201414 39134
rect 200794 3454 201414 38898
rect 200794 3218 200826 3454
rect 201062 3218 201146 3454
rect 201382 3218 201414 3454
rect 200794 3134 201414 3218
rect 200794 2898 200826 3134
rect 201062 2898 201146 3134
rect 201382 2898 201414 3134
rect 200794 -346 201414 2898
rect 200794 -582 200826 -346
rect 201062 -582 201146 -346
rect 201382 -582 201414 -346
rect 200794 -666 201414 -582
rect 200794 -902 200826 -666
rect 201062 -902 201146 -666
rect 201382 -902 201414 -666
rect 200794 -1894 201414 -902
rect 201954 680614 202574 711002
rect 211954 710598 212574 711590
rect 211954 710362 211986 710598
rect 212222 710362 212306 710598
rect 212542 710362 212574 710598
rect 211954 710278 212574 710362
rect 211954 710042 211986 710278
rect 212222 710042 212306 710278
rect 212542 710042 212574 710278
rect 208234 708678 208854 709670
rect 208234 708442 208266 708678
rect 208502 708442 208586 708678
rect 208822 708442 208854 708678
rect 208234 708358 208854 708442
rect 208234 708122 208266 708358
rect 208502 708122 208586 708358
rect 208822 708122 208854 708358
rect 201954 680378 201986 680614
rect 202222 680378 202306 680614
rect 202542 680378 202574 680614
rect 201954 680294 202574 680378
rect 201954 680058 201986 680294
rect 202222 680058 202306 680294
rect 202542 680058 202574 680294
rect 201954 644614 202574 680058
rect 201954 644378 201986 644614
rect 202222 644378 202306 644614
rect 202542 644378 202574 644614
rect 201954 644294 202574 644378
rect 201954 644058 201986 644294
rect 202222 644058 202306 644294
rect 202542 644058 202574 644294
rect 201954 608614 202574 644058
rect 201954 608378 201986 608614
rect 202222 608378 202306 608614
rect 202542 608378 202574 608614
rect 201954 608294 202574 608378
rect 201954 608058 201986 608294
rect 202222 608058 202306 608294
rect 202542 608058 202574 608294
rect 201954 572614 202574 608058
rect 201954 572378 201986 572614
rect 202222 572378 202306 572614
rect 202542 572378 202574 572614
rect 201954 572294 202574 572378
rect 201954 572058 201986 572294
rect 202222 572058 202306 572294
rect 202542 572058 202574 572294
rect 201954 536614 202574 572058
rect 201954 536378 201986 536614
rect 202222 536378 202306 536614
rect 202542 536378 202574 536614
rect 201954 536294 202574 536378
rect 201954 536058 201986 536294
rect 202222 536058 202306 536294
rect 202542 536058 202574 536294
rect 201954 500614 202574 536058
rect 201954 500378 201986 500614
rect 202222 500378 202306 500614
rect 202542 500378 202574 500614
rect 201954 500294 202574 500378
rect 201954 500058 201986 500294
rect 202222 500058 202306 500294
rect 202542 500058 202574 500294
rect 201954 464614 202574 500058
rect 201954 464378 201986 464614
rect 202222 464378 202306 464614
rect 202542 464378 202574 464614
rect 201954 464294 202574 464378
rect 201954 464058 201986 464294
rect 202222 464058 202306 464294
rect 202542 464058 202574 464294
rect 201954 428614 202574 464058
rect 201954 428378 201986 428614
rect 202222 428378 202306 428614
rect 202542 428378 202574 428614
rect 201954 428294 202574 428378
rect 201954 428058 201986 428294
rect 202222 428058 202306 428294
rect 202542 428058 202574 428294
rect 201954 392614 202574 428058
rect 201954 392378 201986 392614
rect 202222 392378 202306 392614
rect 202542 392378 202574 392614
rect 201954 392294 202574 392378
rect 201954 392058 201986 392294
rect 202222 392058 202306 392294
rect 202542 392058 202574 392294
rect 201954 356614 202574 392058
rect 201954 356378 201986 356614
rect 202222 356378 202306 356614
rect 202542 356378 202574 356614
rect 201954 356294 202574 356378
rect 201954 356058 201986 356294
rect 202222 356058 202306 356294
rect 202542 356058 202574 356294
rect 201954 320614 202574 356058
rect 201954 320378 201986 320614
rect 202222 320378 202306 320614
rect 202542 320378 202574 320614
rect 201954 320294 202574 320378
rect 201954 320058 201986 320294
rect 202222 320058 202306 320294
rect 202542 320058 202574 320294
rect 201954 284614 202574 320058
rect 201954 284378 201986 284614
rect 202222 284378 202306 284614
rect 202542 284378 202574 284614
rect 201954 284294 202574 284378
rect 201954 284058 201986 284294
rect 202222 284058 202306 284294
rect 202542 284058 202574 284294
rect 201954 248614 202574 284058
rect 201954 248378 201986 248614
rect 202222 248378 202306 248614
rect 202542 248378 202574 248614
rect 201954 248294 202574 248378
rect 201954 248058 201986 248294
rect 202222 248058 202306 248294
rect 202542 248058 202574 248294
rect 201954 212614 202574 248058
rect 201954 212378 201986 212614
rect 202222 212378 202306 212614
rect 202542 212378 202574 212614
rect 201954 212294 202574 212378
rect 201954 212058 201986 212294
rect 202222 212058 202306 212294
rect 202542 212058 202574 212294
rect 201954 176614 202574 212058
rect 201954 176378 201986 176614
rect 202222 176378 202306 176614
rect 202542 176378 202574 176614
rect 201954 176294 202574 176378
rect 201954 176058 201986 176294
rect 202222 176058 202306 176294
rect 202542 176058 202574 176294
rect 201954 140614 202574 176058
rect 201954 140378 201986 140614
rect 202222 140378 202306 140614
rect 202542 140378 202574 140614
rect 201954 140294 202574 140378
rect 201954 140058 201986 140294
rect 202222 140058 202306 140294
rect 202542 140058 202574 140294
rect 201954 104614 202574 140058
rect 201954 104378 201986 104614
rect 202222 104378 202306 104614
rect 202542 104378 202574 104614
rect 201954 104294 202574 104378
rect 201954 104058 201986 104294
rect 202222 104058 202306 104294
rect 202542 104058 202574 104294
rect 201954 68614 202574 104058
rect 201954 68378 201986 68614
rect 202222 68378 202306 68614
rect 202542 68378 202574 68614
rect 201954 68294 202574 68378
rect 201954 68058 201986 68294
rect 202222 68058 202306 68294
rect 202542 68058 202574 68294
rect 201954 32614 202574 68058
rect 201954 32378 201986 32614
rect 202222 32378 202306 32614
rect 202542 32378 202574 32614
rect 201954 32294 202574 32378
rect 201954 32058 201986 32294
rect 202222 32058 202306 32294
rect 202542 32058 202574 32294
rect 198234 -5382 198266 -5146
rect 198502 -5382 198586 -5146
rect 198822 -5382 198854 -5146
rect 198234 -5466 198854 -5382
rect 198234 -5702 198266 -5466
rect 198502 -5702 198586 -5466
rect 198822 -5702 198854 -5466
rect 198234 -5734 198854 -5702
rect 191954 -6342 191986 -6106
rect 192222 -6342 192306 -6106
rect 192542 -6342 192574 -6106
rect 191954 -6426 192574 -6342
rect 191954 -6662 191986 -6426
rect 192222 -6662 192306 -6426
rect 192542 -6662 192574 -6426
rect 191954 -7654 192574 -6662
rect 201954 -7066 202574 32058
rect 204514 706758 205134 707750
rect 204514 706522 204546 706758
rect 204782 706522 204866 706758
rect 205102 706522 205134 706758
rect 204514 706438 205134 706522
rect 204514 706202 204546 706438
rect 204782 706202 204866 706438
rect 205102 706202 205134 706438
rect 204514 691174 205134 706202
rect 204514 690938 204546 691174
rect 204782 690938 204866 691174
rect 205102 690938 205134 691174
rect 204514 690854 205134 690938
rect 204514 690618 204546 690854
rect 204782 690618 204866 690854
rect 205102 690618 205134 690854
rect 204514 655174 205134 690618
rect 204514 654938 204546 655174
rect 204782 654938 204866 655174
rect 205102 654938 205134 655174
rect 204514 654854 205134 654938
rect 204514 654618 204546 654854
rect 204782 654618 204866 654854
rect 205102 654618 205134 654854
rect 204514 619174 205134 654618
rect 204514 618938 204546 619174
rect 204782 618938 204866 619174
rect 205102 618938 205134 619174
rect 204514 618854 205134 618938
rect 204514 618618 204546 618854
rect 204782 618618 204866 618854
rect 205102 618618 205134 618854
rect 204514 583174 205134 618618
rect 204514 582938 204546 583174
rect 204782 582938 204866 583174
rect 205102 582938 205134 583174
rect 204514 582854 205134 582938
rect 204514 582618 204546 582854
rect 204782 582618 204866 582854
rect 205102 582618 205134 582854
rect 204514 547174 205134 582618
rect 204514 546938 204546 547174
rect 204782 546938 204866 547174
rect 205102 546938 205134 547174
rect 204514 546854 205134 546938
rect 204514 546618 204546 546854
rect 204782 546618 204866 546854
rect 205102 546618 205134 546854
rect 204514 511174 205134 546618
rect 204514 510938 204546 511174
rect 204782 510938 204866 511174
rect 205102 510938 205134 511174
rect 204514 510854 205134 510938
rect 204514 510618 204546 510854
rect 204782 510618 204866 510854
rect 205102 510618 205134 510854
rect 204514 475174 205134 510618
rect 204514 474938 204546 475174
rect 204782 474938 204866 475174
rect 205102 474938 205134 475174
rect 204514 474854 205134 474938
rect 204514 474618 204546 474854
rect 204782 474618 204866 474854
rect 205102 474618 205134 474854
rect 204514 439174 205134 474618
rect 204514 438938 204546 439174
rect 204782 438938 204866 439174
rect 205102 438938 205134 439174
rect 204514 438854 205134 438938
rect 204514 438618 204546 438854
rect 204782 438618 204866 438854
rect 205102 438618 205134 438854
rect 204514 403174 205134 438618
rect 204514 402938 204546 403174
rect 204782 402938 204866 403174
rect 205102 402938 205134 403174
rect 204514 402854 205134 402938
rect 204514 402618 204546 402854
rect 204782 402618 204866 402854
rect 205102 402618 205134 402854
rect 204514 367174 205134 402618
rect 204514 366938 204546 367174
rect 204782 366938 204866 367174
rect 205102 366938 205134 367174
rect 204514 366854 205134 366938
rect 204514 366618 204546 366854
rect 204782 366618 204866 366854
rect 205102 366618 205134 366854
rect 204514 331174 205134 366618
rect 204514 330938 204546 331174
rect 204782 330938 204866 331174
rect 205102 330938 205134 331174
rect 204514 330854 205134 330938
rect 204514 330618 204546 330854
rect 204782 330618 204866 330854
rect 205102 330618 205134 330854
rect 204514 295174 205134 330618
rect 204514 294938 204546 295174
rect 204782 294938 204866 295174
rect 205102 294938 205134 295174
rect 204514 294854 205134 294938
rect 204514 294618 204546 294854
rect 204782 294618 204866 294854
rect 205102 294618 205134 294854
rect 204514 259174 205134 294618
rect 204514 258938 204546 259174
rect 204782 258938 204866 259174
rect 205102 258938 205134 259174
rect 204514 258854 205134 258938
rect 204514 258618 204546 258854
rect 204782 258618 204866 258854
rect 205102 258618 205134 258854
rect 204514 223174 205134 258618
rect 204514 222938 204546 223174
rect 204782 222938 204866 223174
rect 205102 222938 205134 223174
rect 204514 222854 205134 222938
rect 204514 222618 204546 222854
rect 204782 222618 204866 222854
rect 205102 222618 205134 222854
rect 204514 187174 205134 222618
rect 204514 186938 204546 187174
rect 204782 186938 204866 187174
rect 205102 186938 205134 187174
rect 204514 186854 205134 186938
rect 204514 186618 204546 186854
rect 204782 186618 204866 186854
rect 205102 186618 205134 186854
rect 204514 151174 205134 186618
rect 204514 150938 204546 151174
rect 204782 150938 204866 151174
rect 205102 150938 205134 151174
rect 204514 150854 205134 150938
rect 204514 150618 204546 150854
rect 204782 150618 204866 150854
rect 205102 150618 205134 150854
rect 204514 115174 205134 150618
rect 204514 114938 204546 115174
rect 204782 114938 204866 115174
rect 205102 114938 205134 115174
rect 204514 114854 205134 114938
rect 204514 114618 204546 114854
rect 204782 114618 204866 114854
rect 205102 114618 205134 114854
rect 204514 79174 205134 114618
rect 204514 78938 204546 79174
rect 204782 78938 204866 79174
rect 205102 78938 205134 79174
rect 204514 78854 205134 78938
rect 204514 78618 204546 78854
rect 204782 78618 204866 78854
rect 205102 78618 205134 78854
rect 204514 43174 205134 78618
rect 204514 42938 204546 43174
rect 204782 42938 204866 43174
rect 205102 42938 205134 43174
rect 204514 42854 205134 42938
rect 204514 42618 204546 42854
rect 204782 42618 204866 42854
rect 205102 42618 205134 42854
rect 204514 7174 205134 42618
rect 204514 6938 204546 7174
rect 204782 6938 204866 7174
rect 205102 6938 205134 7174
rect 204514 6854 205134 6938
rect 204514 6618 204546 6854
rect 204782 6618 204866 6854
rect 205102 6618 205134 6854
rect 204514 -2266 205134 6618
rect 204514 -2502 204546 -2266
rect 204782 -2502 204866 -2266
rect 205102 -2502 205134 -2266
rect 204514 -2586 205134 -2502
rect 204514 -2822 204546 -2586
rect 204782 -2822 204866 -2586
rect 205102 -2822 205134 -2586
rect 204514 -3814 205134 -2822
rect 208234 694894 208854 708122
rect 208234 694658 208266 694894
rect 208502 694658 208586 694894
rect 208822 694658 208854 694894
rect 208234 694574 208854 694658
rect 208234 694338 208266 694574
rect 208502 694338 208586 694574
rect 208822 694338 208854 694574
rect 208234 658894 208854 694338
rect 208234 658658 208266 658894
rect 208502 658658 208586 658894
rect 208822 658658 208854 658894
rect 208234 658574 208854 658658
rect 208234 658338 208266 658574
rect 208502 658338 208586 658574
rect 208822 658338 208854 658574
rect 208234 622894 208854 658338
rect 208234 622658 208266 622894
rect 208502 622658 208586 622894
rect 208822 622658 208854 622894
rect 208234 622574 208854 622658
rect 208234 622338 208266 622574
rect 208502 622338 208586 622574
rect 208822 622338 208854 622574
rect 208234 586894 208854 622338
rect 208234 586658 208266 586894
rect 208502 586658 208586 586894
rect 208822 586658 208854 586894
rect 208234 586574 208854 586658
rect 208234 586338 208266 586574
rect 208502 586338 208586 586574
rect 208822 586338 208854 586574
rect 208234 550894 208854 586338
rect 208234 550658 208266 550894
rect 208502 550658 208586 550894
rect 208822 550658 208854 550894
rect 208234 550574 208854 550658
rect 208234 550338 208266 550574
rect 208502 550338 208586 550574
rect 208822 550338 208854 550574
rect 208234 514894 208854 550338
rect 208234 514658 208266 514894
rect 208502 514658 208586 514894
rect 208822 514658 208854 514894
rect 208234 514574 208854 514658
rect 208234 514338 208266 514574
rect 208502 514338 208586 514574
rect 208822 514338 208854 514574
rect 208234 478894 208854 514338
rect 208234 478658 208266 478894
rect 208502 478658 208586 478894
rect 208822 478658 208854 478894
rect 208234 478574 208854 478658
rect 208234 478338 208266 478574
rect 208502 478338 208586 478574
rect 208822 478338 208854 478574
rect 208234 442894 208854 478338
rect 208234 442658 208266 442894
rect 208502 442658 208586 442894
rect 208822 442658 208854 442894
rect 208234 442574 208854 442658
rect 208234 442338 208266 442574
rect 208502 442338 208586 442574
rect 208822 442338 208854 442574
rect 208234 406894 208854 442338
rect 208234 406658 208266 406894
rect 208502 406658 208586 406894
rect 208822 406658 208854 406894
rect 208234 406574 208854 406658
rect 208234 406338 208266 406574
rect 208502 406338 208586 406574
rect 208822 406338 208854 406574
rect 208234 370894 208854 406338
rect 208234 370658 208266 370894
rect 208502 370658 208586 370894
rect 208822 370658 208854 370894
rect 208234 370574 208854 370658
rect 208234 370338 208266 370574
rect 208502 370338 208586 370574
rect 208822 370338 208854 370574
rect 208234 334894 208854 370338
rect 208234 334658 208266 334894
rect 208502 334658 208586 334894
rect 208822 334658 208854 334894
rect 208234 334574 208854 334658
rect 208234 334338 208266 334574
rect 208502 334338 208586 334574
rect 208822 334338 208854 334574
rect 208234 298894 208854 334338
rect 208234 298658 208266 298894
rect 208502 298658 208586 298894
rect 208822 298658 208854 298894
rect 208234 298574 208854 298658
rect 208234 298338 208266 298574
rect 208502 298338 208586 298574
rect 208822 298338 208854 298574
rect 208234 262894 208854 298338
rect 208234 262658 208266 262894
rect 208502 262658 208586 262894
rect 208822 262658 208854 262894
rect 208234 262574 208854 262658
rect 208234 262338 208266 262574
rect 208502 262338 208586 262574
rect 208822 262338 208854 262574
rect 208234 226894 208854 262338
rect 208234 226658 208266 226894
rect 208502 226658 208586 226894
rect 208822 226658 208854 226894
rect 208234 226574 208854 226658
rect 208234 226338 208266 226574
rect 208502 226338 208586 226574
rect 208822 226338 208854 226574
rect 208234 190894 208854 226338
rect 208234 190658 208266 190894
rect 208502 190658 208586 190894
rect 208822 190658 208854 190894
rect 208234 190574 208854 190658
rect 208234 190338 208266 190574
rect 208502 190338 208586 190574
rect 208822 190338 208854 190574
rect 208234 154894 208854 190338
rect 208234 154658 208266 154894
rect 208502 154658 208586 154894
rect 208822 154658 208854 154894
rect 208234 154574 208854 154658
rect 208234 154338 208266 154574
rect 208502 154338 208586 154574
rect 208822 154338 208854 154574
rect 208234 118894 208854 154338
rect 208234 118658 208266 118894
rect 208502 118658 208586 118894
rect 208822 118658 208854 118894
rect 208234 118574 208854 118658
rect 208234 118338 208266 118574
rect 208502 118338 208586 118574
rect 208822 118338 208854 118574
rect 208234 82894 208854 118338
rect 208234 82658 208266 82894
rect 208502 82658 208586 82894
rect 208822 82658 208854 82894
rect 208234 82574 208854 82658
rect 208234 82338 208266 82574
rect 208502 82338 208586 82574
rect 208822 82338 208854 82574
rect 208234 46894 208854 82338
rect 208234 46658 208266 46894
rect 208502 46658 208586 46894
rect 208822 46658 208854 46894
rect 208234 46574 208854 46658
rect 208234 46338 208266 46574
rect 208502 46338 208586 46574
rect 208822 46338 208854 46574
rect 208234 10894 208854 46338
rect 208234 10658 208266 10894
rect 208502 10658 208586 10894
rect 208822 10658 208854 10894
rect 208234 10574 208854 10658
rect 208234 10338 208266 10574
rect 208502 10338 208586 10574
rect 208822 10338 208854 10574
rect 208234 -4186 208854 10338
rect 210794 705798 211414 705830
rect 210794 705562 210826 705798
rect 211062 705562 211146 705798
rect 211382 705562 211414 705798
rect 210794 705478 211414 705562
rect 210794 705242 210826 705478
rect 211062 705242 211146 705478
rect 211382 705242 211414 705478
rect 210794 669454 211414 705242
rect 210794 669218 210826 669454
rect 211062 669218 211146 669454
rect 211382 669218 211414 669454
rect 210794 669134 211414 669218
rect 210794 668898 210826 669134
rect 211062 668898 211146 669134
rect 211382 668898 211414 669134
rect 210794 633454 211414 668898
rect 210794 633218 210826 633454
rect 211062 633218 211146 633454
rect 211382 633218 211414 633454
rect 210794 633134 211414 633218
rect 210794 632898 210826 633134
rect 211062 632898 211146 633134
rect 211382 632898 211414 633134
rect 210794 597454 211414 632898
rect 210794 597218 210826 597454
rect 211062 597218 211146 597454
rect 211382 597218 211414 597454
rect 210794 597134 211414 597218
rect 210794 596898 210826 597134
rect 211062 596898 211146 597134
rect 211382 596898 211414 597134
rect 210794 561454 211414 596898
rect 210794 561218 210826 561454
rect 211062 561218 211146 561454
rect 211382 561218 211414 561454
rect 210794 561134 211414 561218
rect 210794 560898 210826 561134
rect 211062 560898 211146 561134
rect 211382 560898 211414 561134
rect 210794 525454 211414 560898
rect 210794 525218 210826 525454
rect 211062 525218 211146 525454
rect 211382 525218 211414 525454
rect 210794 525134 211414 525218
rect 210794 524898 210826 525134
rect 211062 524898 211146 525134
rect 211382 524898 211414 525134
rect 210794 489454 211414 524898
rect 210794 489218 210826 489454
rect 211062 489218 211146 489454
rect 211382 489218 211414 489454
rect 210794 489134 211414 489218
rect 210794 488898 210826 489134
rect 211062 488898 211146 489134
rect 211382 488898 211414 489134
rect 210794 453454 211414 488898
rect 210794 453218 210826 453454
rect 211062 453218 211146 453454
rect 211382 453218 211414 453454
rect 210794 453134 211414 453218
rect 210794 452898 210826 453134
rect 211062 452898 211146 453134
rect 211382 452898 211414 453134
rect 210794 417454 211414 452898
rect 210794 417218 210826 417454
rect 211062 417218 211146 417454
rect 211382 417218 211414 417454
rect 210794 417134 211414 417218
rect 210794 416898 210826 417134
rect 211062 416898 211146 417134
rect 211382 416898 211414 417134
rect 210794 381454 211414 416898
rect 210794 381218 210826 381454
rect 211062 381218 211146 381454
rect 211382 381218 211414 381454
rect 210794 381134 211414 381218
rect 210794 380898 210826 381134
rect 211062 380898 211146 381134
rect 211382 380898 211414 381134
rect 210794 345454 211414 380898
rect 210794 345218 210826 345454
rect 211062 345218 211146 345454
rect 211382 345218 211414 345454
rect 210794 345134 211414 345218
rect 210794 344898 210826 345134
rect 211062 344898 211146 345134
rect 211382 344898 211414 345134
rect 210794 309454 211414 344898
rect 210794 309218 210826 309454
rect 211062 309218 211146 309454
rect 211382 309218 211414 309454
rect 210794 309134 211414 309218
rect 210794 308898 210826 309134
rect 211062 308898 211146 309134
rect 211382 308898 211414 309134
rect 210794 273454 211414 308898
rect 210794 273218 210826 273454
rect 211062 273218 211146 273454
rect 211382 273218 211414 273454
rect 210794 273134 211414 273218
rect 210794 272898 210826 273134
rect 211062 272898 211146 273134
rect 211382 272898 211414 273134
rect 210794 237454 211414 272898
rect 210794 237218 210826 237454
rect 211062 237218 211146 237454
rect 211382 237218 211414 237454
rect 210794 237134 211414 237218
rect 210794 236898 210826 237134
rect 211062 236898 211146 237134
rect 211382 236898 211414 237134
rect 210794 201454 211414 236898
rect 210794 201218 210826 201454
rect 211062 201218 211146 201454
rect 211382 201218 211414 201454
rect 210794 201134 211414 201218
rect 210794 200898 210826 201134
rect 211062 200898 211146 201134
rect 211382 200898 211414 201134
rect 210794 165454 211414 200898
rect 210794 165218 210826 165454
rect 211062 165218 211146 165454
rect 211382 165218 211414 165454
rect 210794 165134 211414 165218
rect 210794 164898 210826 165134
rect 211062 164898 211146 165134
rect 211382 164898 211414 165134
rect 210794 129454 211414 164898
rect 210794 129218 210826 129454
rect 211062 129218 211146 129454
rect 211382 129218 211414 129454
rect 210794 129134 211414 129218
rect 210794 128898 210826 129134
rect 211062 128898 211146 129134
rect 211382 128898 211414 129134
rect 210794 93454 211414 128898
rect 210794 93218 210826 93454
rect 211062 93218 211146 93454
rect 211382 93218 211414 93454
rect 210794 93134 211414 93218
rect 210794 92898 210826 93134
rect 211062 92898 211146 93134
rect 211382 92898 211414 93134
rect 210794 57454 211414 92898
rect 210794 57218 210826 57454
rect 211062 57218 211146 57454
rect 211382 57218 211414 57454
rect 210794 57134 211414 57218
rect 210794 56898 210826 57134
rect 211062 56898 211146 57134
rect 211382 56898 211414 57134
rect 210794 21454 211414 56898
rect 210794 21218 210826 21454
rect 211062 21218 211146 21454
rect 211382 21218 211414 21454
rect 210794 21134 211414 21218
rect 210794 20898 210826 21134
rect 211062 20898 211146 21134
rect 211382 20898 211414 21134
rect 210794 -1306 211414 20898
rect 210794 -1542 210826 -1306
rect 211062 -1542 211146 -1306
rect 211382 -1542 211414 -1306
rect 210794 -1626 211414 -1542
rect 210794 -1862 210826 -1626
rect 211062 -1862 211146 -1626
rect 211382 -1862 211414 -1626
rect 210794 -1894 211414 -1862
rect 211954 698614 212574 710042
rect 221954 711558 222574 711590
rect 221954 711322 221986 711558
rect 222222 711322 222306 711558
rect 222542 711322 222574 711558
rect 221954 711238 222574 711322
rect 221954 711002 221986 711238
rect 222222 711002 222306 711238
rect 222542 711002 222574 711238
rect 218234 709638 218854 709670
rect 218234 709402 218266 709638
rect 218502 709402 218586 709638
rect 218822 709402 218854 709638
rect 218234 709318 218854 709402
rect 218234 709082 218266 709318
rect 218502 709082 218586 709318
rect 218822 709082 218854 709318
rect 211954 698378 211986 698614
rect 212222 698378 212306 698614
rect 212542 698378 212574 698614
rect 211954 698294 212574 698378
rect 211954 698058 211986 698294
rect 212222 698058 212306 698294
rect 212542 698058 212574 698294
rect 211954 662614 212574 698058
rect 211954 662378 211986 662614
rect 212222 662378 212306 662614
rect 212542 662378 212574 662614
rect 211954 662294 212574 662378
rect 211954 662058 211986 662294
rect 212222 662058 212306 662294
rect 212542 662058 212574 662294
rect 211954 626614 212574 662058
rect 211954 626378 211986 626614
rect 212222 626378 212306 626614
rect 212542 626378 212574 626614
rect 211954 626294 212574 626378
rect 211954 626058 211986 626294
rect 212222 626058 212306 626294
rect 212542 626058 212574 626294
rect 211954 590614 212574 626058
rect 211954 590378 211986 590614
rect 212222 590378 212306 590614
rect 212542 590378 212574 590614
rect 211954 590294 212574 590378
rect 211954 590058 211986 590294
rect 212222 590058 212306 590294
rect 212542 590058 212574 590294
rect 211954 554614 212574 590058
rect 211954 554378 211986 554614
rect 212222 554378 212306 554614
rect 212542 554378 212574 554614
rect 211954 554294 212574 554378
rect 211954 554058 211986 554294
rect 212222 554058 212306 554294
rect 212542 554058 212574 554294
rect 211954 518614 212574 554058
rect 211954 518378 211986 518614
rect 212222 518378 212306 518614
rect 212542 518378 212574 518614
rect 211954 518294 212574 518378
rect 211954 518058 211986 518294
rect 212222 518058 212306 518294
rect 212542 518058 212574 518294
rect 211954 482614 212574 518058
rect 211954 482378 211986 482614
rect 212222 482378 212306 482614
rect 212542 482378 212574 482614
rect 211954 482294 212574 482378
rect 211954 482058 211986 482294
rect 212222 482058 212306 482294
rect 212542 482058 212574 482294
rect 211954 446614 212574 482058
rect 211954 446378 211986 446614
rect 212222 446378 212306 446614
rect 212542 446378 212574 446614
rect 211954 446294 212574 446378
rect 211954 446058 211986 446294
rect 212222 446058 212306 446294
rect 212542 446058 212574 446294
rect 211954 410614 212574 446058
rect 211954 410378 211986 410614
rect 212222 410378 212306 410614
rect 212542 410378 212574 410614
rect 211954 410294 212574 410378
rect 211954 410058 211986 410294
rect 212222 410058 212306 410294
rect 212542 410058 212574 410294
rect 211954 374614 212574 410058
rect 211954 374378 211986 374614
rect 212222 374378 212306 374614
rect 212542 374378 212574 374614
rect 211954 374294 212574 374378
rect 211954 374058 211986 374294
rect 212222 374058 212306 374294
rect 212542 374058 212574 374294
rect 211954 338614 212574 374058
rect 211954 338378 211986 338614
rect 212222 338378 212306 338614
rect 212542 338378 212574 338614
rect 211954 338294 212574 338378
rect 211954 338058 211986 338294
rect 212222 338058 212306 338294
rect 212542 338058 212574 338294
rect 211954 302614 212574 338058
rect 211954 302378 211986 302614
rect 212222 302378 212306 302614
rect 212542 302378 212574 302614
rect 211954 302294 212574 302378
rect 211954 302058 211986 302294
rect 212222 302058 212306 302294
rect 212542 302058 212574 302294
rect 211954 266614 212574 302058
rect 211954 266378 211986 266614
rect 212222 266378 212306 266614
rect 212542 266378 212574 266614
rect 211954 266294 212574 266378
rect 211954 266058 211986 266294
rect 212222 266058 212306 266294
rect 212542 266058 212574 266294
rect 211954 230614 212574 266058
rect 211954 230378 211986 230614
rect 212222 230378 212306 230614
rect 212542 230378 212574 230614
rect 211954 230294 212574 230378
rect 211954 230058 211986 230294
rect 212222 230058 212306 230294
rect 212542 230058 212574 230294
rect 211954 194614 212574 230058
rect 211954 194378 211986 194614
rect 212222 194378 212306 194614
rect 212542 194378 212574 194614
rect 211954 194294 212574 194378
rect 211954 194058 211986 194294
rect 212222 194058 212306 194294
rect 212542 194058 212574 194294
rect 211954 158614 212574 194058
rect 211954 158378 211986 158614
rect 212222 158378 212306 158614
rect 212542 158378 212574 158614
rect 211954 158294 212574 158378
rect 211954 158058 211986 158294
rect 212222 158058 212306 158294
rect 212542 158058 212574 158294
rect 211954 122614 212574 158058
rect 211954 122378 211986 122614
rect 212222 122378 212306 122614
rect 212542 122378 212574 122614
rect 211954 122294 212574 122378
rect 211954 122058 211986 122294
rect 212222 122058 212306 122294
rect 212542 122058 212574 122294
rect 211954 86614 212574 122058
rect 211954 86378 211986 86614
rect 212222 86378 212306 86614
rect 212542 86378 212574 86614
rect 211954 86294 212574 86378
rect 211954 86058 211986 86294
rect 212222 86058 212306 86294
rect 212542 86058 212574 86294
rect 211954 50614 212574 86058
rect 211954 50378 211986 50614
rect 212222 50378 212306 50614
rect 212542 50378 212574 50614
rect 211954 50294 212574 50378
rect 211954 50058 211986 50294
rect 212222 50058 212306 50294
rect 212542 50058 212574 50294
rect 211954 14614 212574 50058
rect 211954 14378 211986 14614
rect 212222 14378 212306 14614
rect 212542 14378 212574 14614
rect 211954 14294 212574 14378
rect 211954 14058 211986 14294
rect 212222 14058 212306 14294
rect 212542 14058 212574 14294
rect 208234 -4422 208266 -4186
rect 208502 -4422 208586 -4186
rect 208822 -4422 208854 -4186
rect 208234 -4506 208854 -4422
rect 208234 -4742 208266 -4506
rect 208502 -4742 208586 -4506
rect 208822 -4742 208854 -4506
rect 208234 -5734 208854 -4742
rect 201954 -7302 201986 -7066
rect 202222 -7302 202306 -7066
rect 202542 -7302 202574 -7066
rect 201954 -7386 202574 -7302
rect 201954 -7622 201986 -7386
rect 202222 -7622 202306 -7386
rect 202542 -7622 202574 -7386
rect 201954 -7654 202574 -7622
rect 211954 -6106 212574 14058
rect 214514 707718 215134 707750
rect 214514 707482 214546 707718
rect 214782 707482 214866 707718
rect 215102 707482 215134 707718
rect 214514 707398 215134 707482
rect 214514 707162 214546 707398
rect 214782 707162 214866 707398
rect 215102 707162 215134 707398
rect 214514 673174 215134 707162
rect 214514 672938 214546 673174
rect 214782 672938 214866 673174
rect 215102 672938 215134 673174
rect 214514 672854 215134 672938
rect 214514 672618 214546 672854
rect 214782 672618 214866 672854
rect 215102 672618 215134 672854
rect 214514 637174 215134 672618
rect 214514 636938 214546 637174
rect 214782 636938 214866 637174
rect 215102 636938 215134 637174
rect 214514 636854 215134 636938
rect 214514 636618 214546 636854
rect 214782 636618 214866 636854
rect 215102 636618 215134 636854
rect 214514 601174 215134 636618
rect 214514 600938 214546 601174
rect 214782 600938 214866 601174
rect 215102 600938 215134 601174
rect 214514 600854 215134 600938
rect 214514 600618 214546 600854
rect 214782 600618 214866 600854
rect 215102 600618 215134 600854
rect 214514 565174 215134 600618
rect 214514 564938 214546 565174
rect 214782 564938 214866 565174
rect 215102 564938 215134 565174
rect 214514 564854 215134 564938
rect 214514 564618 214546 564854
rect 214782 564618 214866 564854
rect 215102 564618 215134 564854
rect 214514 529174 215134 564618
rect 214514 528938 214546 529174
rect 214782 528938 214866 529174
rect 215102 528938 215134 529174
rect 214514 528854 215134 528938
rect 214514 528618 214546 528854
rect 214782 528618 214866 528854
rect 215102 528618 215134 528854
rect 214514 493174 215134 528618
rect 214514 492938 214546 493174
rect 214782 492938 214866 493174
rect 215102 492938 215134 493174
rect 214514 492854 215134 492938
rect 214514 492618 214546 492854
rect 214782 492618 214866 492854
rect 215102 492618 215134 492854
rect 214514 457174 215134 492618
rect 214514 456938 214546 457174
rect 214782 456938 214866 457174
rect 215102 456938 215134 457174
rect 214514 456854 215134 456938
rect 214514 456618 214546 456854
rect 214782 456618 214866 456854
rect 215102 456618 215134 456854
rect 214514 421174 215134 456618
rect 214514 420938 214546 421174
rect 214782 420938 214866 421174
rect 215102 420938 215134 421174
rect 214514 420854 215134 420938
rect 214514 420618 214546 420854
rect 214782 420618 214866 420854
rect 215102 420618 215134 420854
rect 214514 385174 215134 420618
rect 214514 384938 214546 385174
rect 214782 384938 214866 385174
rect 215102 384938 215134 385174
rect 214514 384854 215134 384938
rect 214514 384618 214546 384854
rect 214782 384618 214866 384854
rect 215102 384618 215134 384854
rect 214514 349174 215134 384618
rect 214514 348938 214546 349174
rect 214782 348938 214866 349174
rect 215102 348938 215134 349174
rect 214514 348854 215134 348938
rect 214514 348618 214546 348854
rect 214782 348618 214866 348854
rect 215102 348618 215134 348854
rect 214514 313174 215134 348618
rect 214514 312938 214546 313174
rect 214782 312938 214866 313174
rect 215102 312938 215134 313174
rect 214514 312854 215134 312938
rect 214514 312618 214546 312854
rect 214782 312618 214866 312854
rect 215102 312618 215134 312854
rect 214514 277174 215134 312618
rect 214514 276938 214546 277174
rect 214782 276938 214866 277174
rect 215102 276938 215134 277174
rect 214514 276854 215134 276938
rect 214514 276618 214546 276854
rect 214782 276618 214866 276854
rect 215102 276618 215134 276854
rect 214514 241174 215134 276618
rect 214514 240938 214546 241174
rect 214782 240938 214866 241174
rect 215102 240938 215134 241174
rect 214514 240854 215134 240938
rect 214514 240618 214546 240854
rect 214782 240618 214866 240854
rect 215102 240618 215134 240854
rect 214514 205174 215134 240618
rect 214514 204938 214546 205174
rect 214782 204938 214866 205174
rect 215102 204938 215134 205174
rect 214514 204854 215134 204938
rect 214514 204618 214546 204854
rect 214782 204618 214866 204854
rect 215102 204618 215134 204854
rect 214514 169174 215134 204618
rect 214514 168938 214546 169174
rect 214782 168938 214866 169174
rect 215102 168938 215134 169174
rect 214514 168854 215134 168938
rect 214514 168618 214546 168854
rect 214782 168618 214866 168854
rect 215102 168618 215134 168854
rect 214514 133174 215134 168618
rect 214514 132938 214546 133174
rect 214782 132938 214866 133174
rect 215102 132938 215134 133174
rect 214514 132854 215134 132938
rect 214514 132618 214546 132854
rect 214782 132618 214866 132854
rect 215102 132618 215134 132854
rect 214514 97174 215134 132618
rect 214514 96938 214546 97174
rect 214782 96938 214866 97174
rect 215102 96938 215134 97174
rect 214514 96854 215134 96938
rect 214514 96618 214546 96854
rect 214782 96618 214866 96854
rect 215102 96618 215134 96854
rect 214514 61174 215134 96618
rect 214514 60938 214546 61174
rect 214782 60938 214866 61174
rect 215102 60938 215134 61174
rect 214514 60854 215134 60938
rect 214514 60618 214546 60854
rect 214782 60618 214866 60854
rect 215102 60618 215134 60854
rect 214514 25174 215134 60618
rect 214514 24938 214546 25174
rect 214782 24938 214866 25174
rect 215102 24938 215134 25174
rect 214514 24854 215134 24938
rect 214514 24618 214546 24854
rect 214782 24618 214866 24854
rect 215102 24618 215134 24854
rect 214514 -3226 215134 24618
rect 214514 -3462 214546 -3226
rect 214782 -3462 214866 -3226
rect 215102 -3462 215134 -3226
rect 214514 -3546 215134 -3462
rect 214514 -3782 214546 -3546
rect 214782 -3782 214866 -3546
rect 215102 -3782 215134 -3546
rect 214514 -3814 215134 -3782
rect 218234 676894 218854 709082
rect 218234 676658 218266 676894
rect 218502 676658 218586 676894
rect 218822 676658 218854 676894
rect 218234 676574 218854 676658
rect 218234 676338 218266 676574
rect 218502 676338 218586 676574
rect 218822 676338 218854 676574
rect 218234 640894 218854 676338
rect 218234 640658 218266 640894
rect 218502 640658 218586 640894
rect 218822 640658 218854 640894
rect 218234 640574 218854 640658
rect 218234 640338 218266 640574
rect 218502 640338 218586 640574
rect 218822 640338 218854 640574
rect 218234 604894 218854 640338
rect 218234 604658 218266 604894
rect 218502 604658 218586 604894
rect 218822 604658 218854 604894
rect 218234 604574 218854 604658
rect 218234 604338 218266 604574
rect 218502 604338 218586 604574
rect 218822 604338 218854 604574
rect 218234 568894 218854 604338
rect 218234 568658 218266 568894
rect 218502 568658 218586 568894
rect 218822 568658 218854 568894
rect 218234 568574 218854 568658
rect 218234 568338 218266 568574
rect 218502 568338 218586 568574
rect 218822 568338 218854 568574
rect 218234 532894 218854 568338
rect 218234 532658 218266 532894
rect 218502 532658 218586 532894
rect 218822 532658 218854 532894
rect 218234 532574 218854 532658
rect 218234 532338 218266 532574
rect 218502 532338 218586 532574
rect 218822 532338 218854 532574
rect 218234 496894 218854 532338
rect 218234 496658 218266 496894
rect 218502 496658 218586 496894
rect 218822 496658 218854 496894
rect 218234 496574 218854 496658
rect 218234 496338 218266 496574
rect 218502 496338 218586 496574
rect 218822 496338 218854 496574
rect 218234 460894 218854 496338
rect 218234 460658 218266 460894
rect 218502 460658 218586 460894
rect 218822 460658 218854 460894
rect 218234 460574 218854 460658
rect 218234 460338 218266 460574
rect 218502 460338 218586 460574
rect 218822 460338 218854 460574
rect 218234 424894 218854 460338
rect 218234 424658 218266 424894
rect 218502 424658 218586 424894
rect 218822 424658 218854 424894
rect 218234 424574 218854 424658
rect 218234 424338 218266 424574
rect 218502 424338 218586 424574
rect 218822 424338 218854 424574
rect 218234 388894 218854 424338
rect 218234 388658 218266 388894
rect 218502 388658 218586 388894
rect 218822 388658 218854 388894
rect 218234 388574 218854 388658
rect 218234 388338 218266 388574
rect 218502 388338 218586 388574
rect 218822 388338 218854 388574
rect 218234 352894 218854 388338
rect 218234 352658 218266 352894
rect 218502 352658 218586 352894
rect 218822 352658 218854 352894
rect 218234 352574 218854 352658
rect 218234 352338 218266 352574
rect 218502 352338 218586 352574
rect 218822 352338 218854 352574
rect 218234 316894 218854 352338
rect 218234 316658 218266 316894
rect 218502 316658 218586 316894
rect 218822 316658 218854 316894
rect 218234 316574 218854 316658
rect 218234 316338 218266 316574
rect 218502 316338 218586 316574
rect 218822 316338 218854 316574
rect 218234 280894 218854 316338
rect 218234 280658 218266 280894
rect 218502 280658 218586 280894
rect 218822 280658 218854 280894
rect 218234 280574 218854 280658
rect 218234 280338 218266 280574
rect 218502 280338 218586 280574
rect 218822 280338 218854 280574
rect 218234 244894 218854 280338
rect 218234 244658 218266 244894
rect 218502 244658 218586 244894
rect 218822 244658 218854 244894
rect 218234 244574 218854 244658
rect 218234 244338 218266 244574
rect 218502 244338 218586 244574
rect 218822 244338 218854 244574
rect 218234 208894 218854 244338
rect 218234 208658 218266 208894
rect 218502 208658 218586 208894
rect 218822 208658 218854 208894
rect 218234 208574 218854 208658
rect 218234 208338 218266 208574
rect 218502 208338 218586 208574
rect 218822 208338 218854 208574
rect 218234 172894 218854 208338
rect 218234 172658 218266 172894
rect 218502 172658 218586 172894
rect 218822 172658 218854 172894
rect 218234 172574 218854 172658
rect 218234 172338 218266 172574
rect 218502 172338 218586 172574
rect 218822 172338 218854 172574
rect 218234 136894 218854 172338
rect 218234 136658 218266 136894
rect 218502 136658 218586 136894
rect 218822 136658 218854 136894
rect 218234 136574 218854 136658
rect 218234 136338 218266 136574
rect 218502 136338 218586 136574
rect 218822 136338 218854 136574
rect 218234 100894 218854 136338
rect 218234 100658 218266 100894
rect 218502 100658 218586 100894
rect 218822 100658 218854 100894
rect 218234 100574 218854 100658
rect 218234 100338 218266 100574
rect 218502 100338 218586 100574
rect 218822 100338 218854 100574
rect 218234 64894 218854 100338
rect 218234 64658 218266 64894
rect 218502 64658 218586 64894
rect 218822 64658 218854 64894
rect 218234 64574 218854 64658
rect 218234 64338 218266 64574
rect 218502 64338 218586 64574
rect 218822 64338 218854 64574
rect 218234 28894 218854 64338
rect 218234 28658 218266 28894
rect 218502 28658 218586 28894
rect 218822 28658 218854 28894
rect 218234 28574 218854 28658
rect 218234 28338 218266 28574
rect 218502 28338 218586 28574
rect 218822 28338 218854 28574
rect 218234 -5146 218854 28338
rect 220794 704838 221414 705830
rect 220794 704602 220826 704838
rect 221062 704602 221146 704838
rect 221382 704602 221414 704838
rect 220794 704518 221414 704602
rect 220794 704282 220826 704518
rect 221062 704282 221146 704518
rect 221382 704282 221414 704518
rect 220794 687454 221414 704282
rect 220794 687218 220826 687454
rect 221062 687218 221146 687454
rect 221382 687218 221414 687454
rect 220794 687134 221414 687218
rect 220794 686898 220826 687134
rect 221062 686898 221146 687134
rect 221382 686898 221414 687134
rect 220794 651454 221414 686898
rect 220794 651218 220826 651454
rect 221062 651218 221146 651454
rect 221382 651218 221414 651454
rect 220794 651134 221414 651218
rect 220794 650898 220826 651134
rect 221062 650898 221146 651134
rect 221382 650898 221414 651134
rect 220794 615454 221414 650898
rect 220794 615218 220826 615454
rect 221062 615218 221146 615454
rect 221382 615218 221414 615454
rect 220794 615134 221414 615218
rect 220794 614898 220826 615134
rect 221062 614898 221146 615134
rect 221382 614898 221414 615134
rect 220794 579454 221414 614898
rect 220794 579218 220826 579454
rect 221062 579218 221146 579454
rect 221382 579218 221414 579454
rect 220794 579134 221414 579218
rect 220794 578898 220826 579134
rect 221062 578898 221146 579134
rect 221382 578898 221414 579134
rect 220794 543454 221414 578898
rect 220794 543218 220826 543454
rect 221062 543218 221146 543454
rect 221382 543218 221414 543454
rect 220794 543134 221414 543218
rect 220794 542898 220826 543134
rect 221062 542898 221146 543134
rect 221382 542898 221414 543134
rect 220794 507454 221414 542898
rect 220794 507218 220826 507454
rect 221062 507218 221146 507454
rect 221382 507218 221414 507454
rect 220794 507134 221414 507218
rect 220794 506898 220826 507134
rect 221062 506898 221146 507134
rect 221382 506898 221414 507134
rect 220794 471454 221414 506898
rect 220794 471218 220826 471454
rect 221062 471218 221146 471454
rect 221382 471218 221414 471454
rect 220794 471134 221414 471218
rect 220794 470898 220826 471134
rect 221062 470898 221146 471134
rect 221382 470898 221414 471134
rect 220794 435454 221414 470898
rect 220794 435218 220826 435454
rect 221062 435218 221146 435454
rect 221382 435218 221414 435454
rect 220794 435134 221414 435218
rect 220794 434898 220826 435134
rect 221062 434898 221146 435134
rect 221382 434898 221414 435134
rect 220794 399454 221414 434898
rect 220794 399218 220826 399454
rect 221062 399218 221146 399454
rect 221382 399218 221414 399454
rect 220794 399134 221414 399218
rect 220794 398898 220826 399134
rect 221062 398898 221146 399134
rect 221382 398898 221414 399134
rect 220794 363454 221414 398898
rect 220794 363218 220826 363454
rect 221062 363218 221146 363454
rect 221382 363218 221414 363454
rect 220794 363134 221414 363218
rect 220794 362898 220826 363134
rect 221062 362898 221146 363134
rect 221382 362898 221414 363134
rect 220794 327454 221414 362898
rect 220794 327218 220826 327454
rect 221062 327218 221146 327454
rect 221382 327218 221414 327454
rect 220794 327134 221414 327218
rect 220794 326898 220826 327134
rect 221062 326898 221146 327134
rect 221382 326898 221414 327134
rect 220794 291454 221414 326898
rect 220794 291218 220826 291454
rect 221062 291218 221146 291454
rect 221382 291218 221414 291454
rect 220794 291134 221414 291218
rect 220794 290898 220826 291134
rect 221062 290898 221146 291134
rect 221382 290898 221414 291134
rect 220794 255454 221414 290898
rect 220794 255218 220826 255454
rect 221062 255218 221146 255454
rect 221382 255218 221414 255454
rect 220794 255134 221414 255218
rect 220794 254898 220826 255134
rect 221062 254898 221146 255134
rect 221382 254898 221414 255134
rect 220794 219454 221414 254898
rect 220794 219218 220826 219454
rect 221062 219218 221146 219454
rect 221382 219218 221414 219454
rect 220794 219134 221414 219218
rect 220794 218898 220826 219134
rect 221062 218898 221146 219134
rect 221382 218898 221414 219134
rect 220794 183454 221414 218898
rect 220794 183218 220826 183454
rect 221062 183218 221146 183454
rect 221382 183218 221414 183454
rect 220794 183134 221414 183218
rect 220794 182898 220826 183134
rect 221062 182898 221146 183134
rect 221382 182898 221414 183134
rect 220794 147454 221414 182898
rect 220794 147218 220826 147454
rect 221062 147218 221146 147454
rect 221382 147218 221414 147454
rect 220794 147134 221414 147218
rect 220794 146898 220826 147134
rect 221062 146898 221146 147134
rect 221382 146898 221414 147134
rect 220794 111454 221414 146898
rect 220794 111218 220826 111454
rect 221062 111218 221146 111454
rect 221382 111218 221414 111454
rect 220794 111134 221414 111218
rect 220794 110898 220826 111134
rect 221062 110898 221146 111134
rect 221382 110898 221414 111134
rect 220794 75454 221414 110898
rect 220794 75218 220826 75454
rect 221062 75218 221146 75454
rect 221382 75218 221414 75454
rect 220794 75134 221414 75218
rect 220794 74898 220826 75134
rect 221062 74898 221146 75134
rect 221382 74898 221414 75134
rect 220794 39454 221414 74898
rect 220794 39218 220826 39454
rect 221062 39218 221146 39454
rect 221382 39218 221414 39454
rect 220794 39134 221414 39218
rect 220794 38898 220826 39134
rect 221062 38898 221146 39134
rect 221382 38898 221414 39134
rect 220794 3454 221414 38898
rect 220794 3218 220826 3454
rect 221062 3218 221146 3454
rect 221382 3218 221414 3454
rect 220794 3134 221414 3218
rect 220794 2898 220826 3134
rect 221062 2898 221146 3134
rect 221382 2898 221414 3134
rect 220794 -346 221414 2898
rect 220794 -582 220826 -346
rect 221062 -582 221146 -346
rect 221382 -582 221414 -346
rect 220794 -666 221414 -582
rect 220794 -902 220826 -666
rect 221062 -902 221146 -666
rect 221382 -902 221414 -666
rect 220794 -1894 221414 -902
rect 221954 680614 222574 711002
rect 231954 710598 232574 711590
rect 231954 710362 231986 710598
rect 232222 710362 232306 710598
rect 232542 710362 232574 710598
rect 231954 710278 232574 710362
rect 231954 710042 231986 710278
rect 232222 710042 232306 710278
rect 232542 710042 232574 710278
rect 228234 708678 228854 709670
rect 228234 708442 228266 708678
rect 228502 708442 228586 708678
rect 228822 708442 228854 708678
rect 228234 708358 228854 708442
rect 228234 708122 228266 708358
rect 228502 708122 228586 708358
rect 228822 708122 228854 708358
rect 221954 680378 221986 680614
rect 222222 680378 222306 680614
rect 222542 680378 222574 680614
rect 221954 680294 222574 680378
rect 221954 680058 221986 680294
rect 222222 680058 222306 680294
rect 222542 680058 222574 680294
rect 221954 644614 222574 680058
rect 221954 644378 221986 644614
rect 222222 644378 222306 644614
rect 222542 644378 222574 644614
rect 221954 644294 222574 644378
rect 221954 644058 221986 644294
rect 222222 644058 222306 644294
rect 222542 644058 222574 644294
rect 221954 608614 222574 644058
rect 221954 608378 221986 608614
rect 222222 608378 222306 608614
rect 222542 608378 222574 608614
rect 221954 608294 222574 608378
rect 221954 608058 221986 608294
rect 222222 608058 222306 608294
rect 222542 608058 222574 608294
rect 221954 572614 222574 608058
rect 221954 572378 221986 572614
rect 222222 572378 222306 572614
rect 222542 572378 222574 572614
rect 221954 572294 222574 572378
rect 221954 572058 221986 572294
rect 222222 572058 222306 572294
rect 222542 572058 222574 572294
rect 221954 536614 222574 572058
rect 221954 536378 221986 536614
rect 222222 536378 222306 536614
rect 222542 536378 222574 536614
rect 221954 536294 222574 536378
rect 221954 536058 221986 536294
rect 222222 536058 222306 536294
rect 222542 536058 222574 536294
rect 221954 500614 222574 536058
rect 221954 500378 221986 500614
rect 222222 500378 222306 500614
rect 222542 500378 222574 500614
rect 221954 500294 222574 500378
rect 221954 500058 221986 500294
rect 222222 500058 222306 500294
rect 222542 500058 222574 500294
rect 221954 464614 222574 500058
rect 221954 464378 221986 464614
rect 222222 464378 222306 464614
rect 222542 464378 222574 464614
rect 221954 464294 222574 464378
rect 221954 464058 221986 464294
rect 222222 464058 222306 464294
rect 222542 464058 222574 464294
rect 221954 428614 222574 464058
rect 221954 428378 221986 428614
rect 222222 428378 222306 428614
rect 222542 428378 222574 428614
rect 221954 428294 222574 428378
rect 221954 428058 221986 428294
rect 222222 428058 222306 428294
rect 222542 428058 222574 428294
rect 221954 392614 222574 428058
rect 221954 392378 221986 392614
rect 222222 392378 222306 392614
rect 222542 392378 222574 392614
rect 221954 392294 222574 392378
rect 221954 392058 221986 392294
rect 222222 392058 222306 392294
rect 222542 392058 222574 392294
rect 221954 356614 222574 392058
rect 221954 356378 221986 356614
rect 222222 356378 222306 356614
rect 222542 356378 222574 356614
rect 221954 356294 222574 356378
rect 221954 356058 221986 356294
rect 222222 356058 222306 356294
rect 222542 356058 222574 356294
rect 221954 320614 222574 356058
rect 221954 320378 221986 320614
rect 222222 320378 222306 320614
rect 222542 320378 222574 320614
rect 221954 320294 222574 320378
rect 221954 320058 221986 320294
rect 222222 320058 222306 320294
rect 222542 320058 222574 320294
rect 221954 284614 222574 320058
rect 221954 284378 221986 284614
rect 222222 284378 222306 284614
rect 222542 284378 222574 284614
rect 221954 284294 222574 284378
rect 221954 284058 221986 284294
rect 222222 284058 222306 284294
rect 222542 284058 222574 284294
rect 221954 248614 222574 284058
rect 221954 248378 221986 248614
rect 222222 248378 222306 248614
rect 222542 248378 222574 248614
rect 221954 248294 222574 248378
rect 221954 248058 221986 248294
rect 222222 248058 222306 248294
rect 222542 248058 222574 248294
rect 221954 212614 222574 248058
rect 221954 212378 221986 212614
rect 222222 212378 222306 212614
rect 222542 212378 222574 212614
rect 221954 212294 222574 212378
rect 221954 212058 221986 212294
rect 222222 212058 222306 212294
rect 222542 212058 222574 212294
rect 221954 176614 222574 212058
rect 221954 176378 221986 176614
rect 222222 176378 222306 176614
rect 222542 176378 222574 176614
rect 221954 176294 222574 176378
rect 221954 176058 221986 176294
rect 222222 176058 222306 176294
rect 222542 176058 222574 176294
rect 221954 140614 222574 176058
rect 221954 140378 221986 140614
rect 222222 140378 222306 140614
rect 222542 140378 222574 140614
rect 221954 140294 222574 140378
rect 221954 140058 221986 140294
rect 222222 140058 222306 140294
rect 222542 140058 222574 140294
rect 221954 104614 222574 140058
rect 221954 104378 221986 104614
rect 222222 104378 222306 104614
rect 222542 104378 222574 104614
rect 221954 104294 222574 104378
rect 221954 104058 221986 104294
rect 222222 104058 222306 104294
rect 222542 104058 222574 104294
rect 221954 68614 222574 104058
rect 221954 68378 221986 68614
rect 222222 68378 222306 68614
rect 222542 68378 222574 68614
rect 221954 68294 222574 68378
rect 221954 68058 221986 68294
rect 222222 68058 222306 68294
rect 222542 68058 222574 68294
rect 221954 32614 222574 68058
rect 221954 32378 221986 32614
rect 222222 32378 222306 32614
rect 222542 32378 222574 32614
rect 221954 32294 222574 32378
rect 221954 32058 221986 32294
rect 222222 32058 222306 32294
rect 222542 32058 222574 32294
rect 218234 -5382 218266 -5146
rect 218502 -5382 218586 -5146
rect 218822 -5382 218854 -5146
rect 218234 -5466 218854 -5382
rect 218234 -5702 218266 -5466
rect 218502 -5702 218586 -5466
rect 218822 -5702 218854 -5466
rect 218234 -5734 218854 -5702
rect 211954 -6342 211986 -6106
rect 212222 -6342 212306 -6106
rect 212542 -6342 212574 -6106
rect 211954 -6426 212574 -6342
rect 211954 -6662 211986 -6426
rect 212222 -6662 212306 -6426
rect 212542 -6662 212574 -6426
rect 211954 -7654 212574 -6662
rect 221954 -7066 222574 32058
rect 224514 706758 225134 707750
rect 224514 706522 224546 706758
rect 224782 706522 224866 706758
rect 225102 706522 225134 706758
rect 224514 706438 225134 706522
rect 224514 706202 224546 706438
rect 224782 706202 224866 706438
rect 225102 706202 225134 706438
rect 224514 691174 225134 706202
rect 224514 690938 224546 691174
rect 224782 690938 224866 691174
rect 225102 690938 225134 691174
rect 224514 690854 225134 690938
rect 224514 690618 224546 690854
rect 224782 690618 224866 690854
rect 225102 690618 225134 690854
rect 224514 655174 225134 690618
rect 224514 654938 224546 655174
rect 224782 654938 224866 655174
rect 225102 654938 225134 655174
rect 224514 654854 225134 654938
rect 224514 654618 224546 654854
rect 224782 654618 224866 654854
rect 225102 654618 225134 654854
rect 224514 619174 225134 654618
rect 224514 618938 224546 619174
rect 224782 618938 224866 619174
rect 225102 618938 225134 619174
rect 224514 618854 225134 618938
rect 224514 618618 224546 618854
rect 224782 618618 224866 618854
rect 225102 618618 225134 618854
rect 224514 583174 225134 618618
rect 224514 582938 224546 583174
rect 224782 582938 224866 583174
rect 225102 582938 225134 583174
rect 224514 582854 225134 582938
rect 224514 582618 224546 582854
rect 224782 582618 224866 582854
rect 225102 582618 225134 582854
rect 224514 547174 225134 582618
rect 224514 546938 224546 547174
rect 224782 546938 224866 547174
rect 225102 546938 225134 547174
rect 224514 546854 225134 546938
rect 224514 546618 224546 546854
rect 224782 546618 224866 546854
rect 225102 546618 225134 546854
rect 224514 511174 225134 546618
rect 224514 510938 224546 511174
rect 224782 510938 224866 511174
rect 225102 510938 225134 511174
rect 224514 510854 225134 510938
rect 224514 510618 224546 510854
rect 224782 510618 224866 510854
rect 225102 510618 225134 510854
rect 224514 475174 225134 510618
rect 224514 474938 224546 475174
rect 224782 474938 224866 475174
rect 225102 474938 225134 475174
rect 224514 474854 225134 474938
rect 224514 474618 224546 474854
rect 224782 474618 224866 474854
rect 225102 474618 225134 474854
rect 224514 439174 225134 474618
rect 224514 438938 224546 439174
rect 224782 438938 224866 439174
rect 225102 438938 225134 439174
rect 224514 438854 225134 438938
rect 224514 438618 224546 438854
rect 224782 438618 224866 438854
rect 225102 438618 225134 438854
rect 224514 403174 225134 438618
rect 224514 402938 224546 403174
rect 224782 402938 224866 403174
rect 225102 402938 225134 403174
rect 224514 402854 225134 402938
rect 224514 402618 224546 402854
rect 224782 402618 224866 402854
rect 225102 402618 225134 402854
rect 224514 367174 225134 402618
rect 224514 366938 224546 367174
rect 224782 366938 224866 367174
rect 225102 366938 225134 367174
rect 224514 366854 225134 366938
rect 224514 366618 224546 366854
rect 224782 366618 224866 366854
rect 225102 366618 225134 366854
rect 224514 331174 225134 366618
rect 224514 330938 224546 331174
rect 224782 330938 224866 331174
rect 225102 330938 225134 331174
rect 224514 330854 225134 330938
rect 224514 330618 224546 330854
rect 224782 330618 224866 330854
rect 225102 330618 225134 330854
rect 224514 295174 225134 330618
rect 224514 294938 224546 295174
rect 224782 294938 224866 295174
rect 225102 294938 225134 295174
rect 224514 294854 225134 294938
rect 224514 294618 224546 294854
rect 224782 294618 224866 294854
rect 225102 294618 225134 294854
rect 224514 259174 225134 294618
rect 224514 258938 224546 259174
rect 224782 258938 224866 259174
rect 225102 258938 225134 259174
rect 224514 258854 225134 258938
rect 224514 258618 224546 258854
rect 224782 258618 224866 258854
rect 225102 258618 225134 258854
rect 224514 223174 225134 258618
rect 224514 222938 224546 223174
rect 224782 222938 224866 223174
rect 225102 222938 225134 223174
rect 224514 222854 225134 222938
rect 224514 222618 224546 222854
rect 224782 222618 224866 222854
rect 225102 222618 225134 222854
rect 224514 187174 225134 222618
rect 224514 186938 224546 187174
rect 224782 186938 224866 187174
rect 225102 186938 225134 187174
rect 224514 186854 225134 186938
rect 224514 186618 224546 186854
rect 224782 186618 224866 186854
rect 225102 186618 225134 186854
rect 224514 151174 225134 186618
rect 224514 150938 224546 151174
rect 224782 150938 224866 151174
rect 225102 150938 225134 151174
rect 224514 150854 225134 150938
rect 224514 150618 224546 150854
rect 224782 150618 224866 150854
rect 225102 150618 225134 150854
rect 224514 115174 225134 150618
rect 224514 114938 224546 115174
rect 224782 114938 224866 115174
rect 225102 114938 225134 115174
rect 224514 114854 225134 114938
rect 224514 114618 224546 114854
rect 224782 114618 224866 114854
rect 225102 114618 225134 114854
rect 224514 79174 225134 114618
rect 224514 78938 224546 79174
rect 224782 78938 224866 79174
rect 225102 78938 225134 79174
rect 224514 78854 225134 78938
rect 224514 78618 224546 78854
rect 224782 78618 224866 78854
rect 225102 78618 225134 78854
rect 224514 43174 225134 78618
rect 224514 42938 224546 43174
rect 224782 42938 224866 43174
rect 225102 42938 225134 43174
rect 224514 42854 225134 42938
rect 224514 42618 224546 42854
rect 224782 42618 224866 42854
rect 225102 42618 225134 42854
rect 224514 7174 225134 42618
rect 224514 6938 224546 7174
rect 224782 6938 224866 7174
rect 225102 6938 225134 7174
rect 224514 6854 225134 6938
rect 224514 6618 224546 6854
rect 224782 6618 224866 6854
rect 225102 6618 225134 6854
rect 224514 -2266 225134 6618
rect 224514 -2502 224546 -2266
rect 224782 -2502 224866 -2266
rect 225102 -2502 225134 -2266
rect 224514 -2586 225134 -2502
rect 224514 -2822 224546 -2586
rect 224782 -2822 224866 -2586
rect 225102 -2822 225134 -2586
rect 224514 -3814 225134 -2822
rect 228234 694894 228854 708122
rect 228234 694658 228266 694894
rect 228502 694658 228586 694894
rect 228822 694658 228854 694894
rect 228234 694574 228854 694658
rect 228234 694338 228266 694574
rect 228502 694338 228586 694574
rect 228822 694338 228854 694574
rect 228234 658894 228854 694338
rect 228234 658658 228266 658894
rect 228502 658658 228586 658894
rect 228822 658658 228854 658894
rect 228234 658574 228854 658658
rect 228234 658338 228266 658574
rect 228502 658338 228586 658574
rect 228822 658338 228854 658574
rect 228234 622894 228854 658338
rect 228234 622658 228266 622894
rect 228502 622658 228586 622894
rect 228822 622658 228854 622894
rect 228234 622574 228854 622658
rect 228234 622338 228266 622574
rect 228502 622338 228586 622574
rect 228822 622338 228854 622574
rect 228234 586894 228854 622338
rect 228234 586658 228266 586894
rect 228502 586658 228586 586894
rect 228822 586658 228854 586894
rect 228234 586574 228854 586658
rect 228234 586338 228266 586574
rect 228502 586338 228586 586574
rect 228822 586338 228854 586574
rect 228234 550894 228854 586338
rect 228234 550658 228266 550894
rect 228502 550658 228586 550894
rect 228822 550658 228854 550894
rect 228234 550574 228854 550658
rect 228234 550338 228266 550574
rect 228502 550338 228586 550574
rect 228822 550338 228854 550574
rect 228234 514894 228854 550338
rect 228234 514658 228266 514894
rect 228502 514658 228586 514894
rect 228822 514658 228854 514894
rect 228234 514574 228854 514658
rect 228234 514338 228266 514574
rect 228502 514338 228586 514574
rect 228822 514338 228854 514574
rect 228234 478894 228854 514338
rect 228234 478658 228266 478894
rect 228502 478658 228586 478894
rect 228822 478658 228854 478894
rect 228234 478574 228854 478658
rect 228234 478338 228266 478574
rect 228502 478338 228586 478574
rect 228822 478338 228854 478574
rect 228234 442894 228854 478338
rect 228234 442658 228266 442894
rect 228502 442658 228586 442894
rect 228822 442658 228854 442894
rect 228234 442574 228854 442658
rect 228234 442338 228266 442574
rect 228502 442338 228586 442574
rect 228822 442338 228854 442574
rect 228234 406894 228854 442338
rect 228234 406658 228266 406894
rect 228502 406658 228586 406894
rect 228822 406658 228854 406894
rect 228234 406574 228854 406658
rect 228234 406338 228266 406574
rect 228502 406338 228586 406574
rect 228822 406338 228854 406574
rect 228234 370894 228854 406338
rect 228234 370658 228266 370894
rect 228502 370658 228586 370894
rect 228822 370658 228854 370894
rect 228234 370574 228854 370658
rect 228234 370338 228266 370574
rect 228502 370338 228586 370574
rect 228822 370338 228854 370574
rect 228234 334894 228854 370338
rect 228234 334658 228266 334894
rect 228502 334658 228586 334894
rect 228822 334658 228854 334894
rect 228234 334574 228854 334658
rect 228234 334338 228266 334574
rect 228502 334338 228586 334574
rect 228822 334338 228854 334574
rect 228234 298894 228854 334338
rect 228234 298658 228266 298894
rect 228502 298658 228586 298894
rect 228822 298658 228854 298894
rect 228234 298574 228854 298658
rect 228234 298338 228266 298574
rect 228502 298338 228586 298574
rect 228822 298338 228854 298574
rect 228234 262894 228854 298338
rect 228234 262658 228266 262894
rect 228502 262658 228586 262894
rect 228822 262658 228854 262894
rect 228234 262574 228854 262658
rect 228234 262338 228266 262574
rect 228502 262338 228586 262574
rect 228822 262338 228854 262574
rect 228234 226894 228854 262338
rect 228234 226658 228266 226894
rect 228502 226658 228586 226894
rect 228822 226658 228854 226894
rect 228234 226574 228854 226658
rect 228234 226338 228266 226574
rect 228502 226338 228586 226574
rect 228822 226338 228854 226574
rect 228234 190894 228854 226338
rect 228234 190658 228266 190894
rect 228502 190658 228586 190894
rect 228822 190658 228854 190894
rect 228234 190574 228854 190658
rect 228234 190338 228266 190574
rect 228502 190338 228586 190574
rect 228822 190338 228854 190574
rect 228234 154894 228854 190338
rect 228234 154658 228266 154894
rect 228502 154658 228586 154894
rect 228822 154658 228854 154894
rect 228234 154574 228854 154658
rect 228234 154338 228266 154574
rect 228502 154338 228586 154574
rect 228822 154338 228854 154574
rect 228234 118894 228854 154338
rect 228234 118658 228266 118894
rect 228502 118658 228586 118894
rect 228822 118658 228854 118894
rect 228234 118574 228854 118658
rect 228234 118338 228266 118574
rect 228502 118338 228586 118574
rect 228822 118338 228854 118574
rect 228234 82894 228854 118338
rect 228234 82658 228266 82894
rect 228502 82658 228586 82894
rect 228822 82658 228854 82894
rect 228234 82574 228854 82658
rect 228234 82338 228266 82574
rect 228502 82338 228586 82574
rect 228822 82338 228854 82574
rect 228234 46894 228854 82338
rect 228234 46658 228266 46894
rect 228502 46658 228586 46894
rect 228822 46658 228854 46894
rect 228234 46574 228854 46658
rect 228234 46338 228266 46574
rect 228502 46338 228586 46574
rect 228822 46338 228854 46574
rect 228234 10894 228854 46338
rect 228234 10658 228266 10894
rect 228502 10658 228586 10894
rect 228822 10658 228854 10894
rect 228234 10574 228854 10658
rect 228234 10338 228266 10574
rect 228502 10338 228586 10574
rect 228822 10338 228854 10574
rect 228234 -4186 228854 10338
rect 230794 705798 231414 705830
rect 230794 705562 230826 705798
rect 231062 705562 231146 705798
rect 231382 705562 231414 705798
rect 230794 705478 231414 705562
rect 230794 705242 230826 705478
rect 231062 705242 231146 705478
rect 231382 705242 231414 705478
rect 230794 669454 231414 705242
rect 230794 669218 230826 669454
rect 231062 669218 231146 669454
rect 231382 669218 231414 669454
rect 230794 669134 231414 669218
rect 230794 668898 230826 669134
rect 231062 668898 231146 669134
rect 231382 668898 231414 669134
rect 230794 633454 231414 668898
rect 230794 633218 230826 633454
rect 231062 633218 231146 633454
rect 231382 633218 231414 633454
rect 230794 633134 231414 633218
rect 230794 632898 230826 633134
rect 231062 632898 231146 633134
rect 231382 632898 231414 633134
rect 230794 597454 231414 632898
rect 230794 597218 230826 597454
rect 231062 597218 231146 597454
rect 231382 597218 231414 597454
rect 230794 597134 231414 597218
rect 230794 596898 230826 597134
rect 231062 596898 231146 597134
rect 231382 596898 231414 597134
rect 230794 561454 231414 596898
rect 230794 561218 230826 561454
rect 231062 561218 231146 561454
rect 231382 561218 231414 561454
rect 230794 561134 231414 561218
rect 230794 560898 230826 561134
rect 231062 560898 231146 561134
rect 231382 560898 231414 561134
rect 230794 525454 231414 560898
rect 230794 525218 230826 525454
rect 231062 525218 231146 525454
rect 231382 525218 231414 525454
rect 230794 525134 231414 525218
rect 230794 524898 230826 525134
rect 231062 524898 231146 525134
rect 231382 524898 231414 525134
rect 230794 489454 231414 524898
rect 230794 489218 230826 489454
rect 231062 489218 231146 489454
rect 231382 489218 231414 489454
rect 230794 489134 231414 489218
rect 230794 488898 230826 489134
rect 231062 488898 231146 489134
rect 231382 488898 231414 489134
rect 230794 453454 231414 488898
rect 230794 453218 230826 453454
rect 231062 453218 231146 453454
rect 231382 453218 231414 453454
rect 230794 453134 231414 453218
rect 230794 452898 230826 453134
rect 231062 452898 231146 453134
rect 231382 452898 231414 453134
rect 230794 417454 231414 452898
rect 230794 417218 230826 417454
rect 231062 417218 231146 417454
rect 231382 417218 231414 417454
rect 230794 417134 231414 417218
rect 230794 416898 230826 417134
rect 231062 416898 231146 417134
rect 231382 416898 231414 417134
rect 230794 381454 231414 416898
rect 230794 381218 230826 381454
rect 231062 381218 231146 381454
rect 231382 381218 231414 381454
rect 230794 381134 231414 381218
rect 230794 380898 230826 381134
rect 231062 380898 231146 381134
rect 231382 380898 231414 381134
rect 230794 345454 231414 380898
rect 230794 345218 230826 345454
rect 231062 345218 231146 345454
rect 231382 345218 231414 345454
rect 230794 345134 231414 345218
rect 230794 344898 230826 345134
rect 231062 344898 231146 345134
rect 231382 344898 231414 345134
rect 230794 309454 231414 344898
rect 230794 309218 230826 309454
rect 231062 309218 231146 309454
rect 231382 309218 231414 309454
rect 230794 309134 231414 309218
rect 230794 308898 230826 309134
rect 231062 308898 231146 309134
rect 231382 308898 231414 309134
rect 230794 273454 231414 308898
rect 230794 273218 230826 273454
rect 231062 273218 231146 273454
rect 231382 273218 231414 273454
rect 230794 273134 231414 273218
rect 230794 272898 230826 273134
rect 231062 272898 231146 273134
rect 231382 272898 231414 273134
rect 230794 237454 231414 272898
rect 230794 237218 230826 237454
rect 231062 237218 231146 237454
rect 231382 237218 231414 237454
rect 230794 237134 231414 237218
rect 230794 236898 230826 237134
rect 231062 236898 231146 237134
rect 231382 236898 231414 237134
rect 230794 201454 231414 236898
rect 230794 201218 230826 201454
rect 231062 201218 231146 201454
rect 231382 201218 231414 201454
rect 230794 201134 231414 201218
rect 230794 200898 230826 201134
rect 231062 200898 231146 201134
rect 231382 200898 231414 201134
rect 230794 165454 231414 200898
rect 230794 165218 230826 165454
rect 231062 165218 231146 165454
rect 231382 165218 231414 165454
rect 230794 165134 231414 165218
rect 230794 164898 230826 165134
rect 231062 164898 231146 165134
rect 231382 164898 231414 165134
rect 230794 129454 231414 164898
rect 230794 129218 230826 129454
rect 231062 129218 231146 129454
rect 231382 129218 231414 129454
rect 230794 129134 231414 129218
rect 230794 128898 230826 129134
rect 231062 128898 231146 129134
rect 231382 128898 231414 129134
rect 230794 93454 231414 128898
rect 230794 93218 230826 93454
rect 231062 93218 231146 93454
rect 231382 93218 231414 93454
rect 230794 93134 231414 93218
rect 230794 92898 230826 93134
rect 231062 92898 231146 93134
rect 231382 92898 231414 93134
rect 230794 57454 231414 92898
rect 230794 57218 230826 57454
rect 231062 57218 231146 57454
rect 231382 57218 231414 57454
rect 230794 57134 231414 57218
rect 230794 56898 230826 57134
rect 231062 56898 231146 57134
rect 231382 56898 231414 57134
rect 230794 21454 231414 56898
rect 230794 21218 230826 21454
rect 231062 21218 231146 21454
rect 231382 21218 231414 21454
rect 230794 21134 231414 21218
rect 230794 20898 230826 21134
rect 231062 20898 231146 21134
rect 231382 20898 231414 21134
rect 230794 -1306 231414 20898
rect 230794 -1542 230826 -1306
rect 231062 -1542 231146 -1306
rect 231382 -1542 231414 -1306
rect 230794 -1626 231414 -1542
rect 230794 -1862 230826 -1626
rect 231062 -1862 231146 -1626
rect 231382 -1862 231414 -1626
rect 230794 -1894 231414 -1862
rect 231954 698614 232574 710042
rect 241954 711558 242574 711590
rect 241954 711322 241986 711558
rect 242222 711322 242306 711558
rect 242542 711322 242574 711558
rect 241954 711238 242574 711322
rect 241954 711002 241986 711238
rect 242222 711002 242306 711238
rect 242542 711002 242574 711238
rect 238234 709638 238854 709670
rect 238234 709402 238266 709638
rect 238502 709402 238586 709638
rect 238822 709402 238854 709638
rect 238234 709318 238854 709402
rect 238234 709082 238266 709318
rect 238502 709082 238586 709318
rect 238822 709082 238854 709318
rect 231954 698378 231986 698614
rect 232222 698378 232306 698614
rect 232542 698378 232574 698614
rect 231954 698294 232574 698378
rect 231954 698058 231986 698294
rect 232222 698058 232306 698294
rect 232542 698058 232574 698294
rect 231954 662614 232574 698058
rect 231954 662378 231986 662614
rect 232222 662378 232306 662614
rect 232542 662378 232574 662614
rect 231954 662294 232574 662378
rect 231954 662058 231986 662294
rect 232222 662058 232306 662294
rect 232542 662058 232574 662294
rect 231954 626614 232574 662058
rect 231954 626378 231986 626614
rect 232222 626378 232306 626614
rect 232542 626378 232574 626614
rect 231954 626294 232574 626378
rect 231954 626058 231986 626294
rect 232222 626058 232306 626294
rect 232542 626058 232574 626294
rect 231954 590614 232574 626058
rect 231954 590378 231986 590614
rect 232222 590378 232306 590614
rect 232542 590378 232574 590614
rect 231954 590294 232574 590378
rect 231954 590058 231986 590294
rect 232222 590058 232306 590294
rect 232542 590058 232574 590294
rect 231954 554614 232574 590058
rect 231954 554378 231986 554614
rect 232222 554378 232306 554614
rect 232542 554378 232574 554614
rect 231954 554294 232574 554378
rect 231954 554058 231986 554294
rect 232222 554058 232306 554294
rect 232542 554058 232574 554294
rect 231954 518614 232574 554058
rect 231954 518378 231986 518614
rect 232222 518378 232306 518614
rect 232542 518378 232574 518614
rect 231954 518294 232574 518378
rect 231954 518058 231986 518294
rect 232222 518058 232306 518294
rect 232542 518058 232574 518294
rect 231954 482614 232574 518058
rect 231954 482378 231986 482614
rect 232222 482378 232306 482614
rect 232542 482378 232574 482614
rect 231954 482294 232574 482378
rect 231954 482058 231986 482294
rect 232222 482058 232306 482294
rect 232542 482058 232574 482294
rect 231954 446614 232574 482058
rect 231954 446378 231986 446614
rect 232222 446378 232306 446614
rect 232542 446378 232574 446614
rect 231954 446294 232574 446378
rect 231954 446058 231986 446294
rect 232222 446058 232306 446294
rect 232542 446058 232574 446294
rect 231954 410614 232574 446058
rect 231954 410378 231986 410614
rect 232222 410378 232306 410614
rect 232542 410378 232574 410614
rect 231954 410294 232574 410378
rect 231954 410058 231986 410294
rect 232222 410058 232306 410294
rect 232542 410058 232574 410294
rect 231954 374614 232574 410058
rect 231954 374378 231986 374614
rect 232222 374378 232306 374614
rect 232542 374378 232574 374614
rect 231954 374294 232574 374378
rect 231954 374058 231986 374294
rect 232222 374058 232306 374294
rect 232542 374058 232574 374294
rect 231954 338614 232574 374058
rect 231954 338378 231986 338614
rect 232222 338378 232306 338614
rect 232542 338378 232574 338614
rect 231954 338294 232574 338378
rect 231954 338058 231986 338294
rect 232222 338058 232306 338294
rect 232542 338058 232574 338294
rect 231954 302614 232574 338058
rect 231954 302378 231986 302614
rect 232222 302378 232306 302614
rect 232542 302378 232574 302614
rect 231954 302294 232574 302378
rect 231954 302058 231986 302294
rect 232222 302058 232306 302294
rect 232542 302058 232574 302294
rect 231954 266614 232574 302058
rect 231954 266378 231986 266614
rect 232222 266378 232306 266614
rect 232542 266378 232574 266614
rect 231954 266294 232574 266378
rect 231954 266058 231986 266294
rect 232222 266058 232306 266294
rect 232542 266058 232574 266294
rect 231954 230614 232574 266058
rect 231954 230378 231986 230614
rect 232222 230378 232306 230614
rect 232542 230378 232574 230614
rect 231954 230294 232574 230378
rect 231954 230058 231986 230294
rect 232222 230058 232306 230294
rect 232542 230058 232574 230294
rect 231954 194614 232574 230058
rect 231954 194378 231986 194614
rect 232222 194378 232306 194614
rect 232542 194378 232574 194614
rect 231954 194294 232574 194378
rect 231954 194058 231986 194294
rect 232222 194058 232306 194294
rect 232542 194058 232574 194294
rect 231954 158614 232574 194058
rect 231954 158378 231986 158614
rect 232222 158378 232306 158614
rect 232542 158378 232574 158614
rect 231954 158294 232574 158378
rect 231954 158058 231986 158294
rect 232222 158058 232306 158294
rect 232542 158058 232574 158294
rect 231954 122614 232574 158058
rect 231954 122378 231986 122614
rect 232222 122378 232306 122614
rect 232542 122378 232574 122614
rect 231954 122294 232574 122378
rect 231954 122058 231986 122294
rect 232222 122058 232306 122294
rect 232542 122058 232574 122294
rect 231954 86614 232574 122058
rect 231954 86378 231986 86614
rect 232222 86378 232306 86614
rect 232542 86378 232574 86614
rect 231954 86294 232574 86378
rect 231954 86058 231986 86294
rect 232222 86058 232306 86294
rect 232542 86058 232574 86294
rect 231954 50614 232574 86058
rect 231954 50378 231986 50614
rect 232222 50378 232306 50614
rect 232542 50378 232574 50614
rect 231954 50294 232574 50378
rect 231954 50058 231986 50294
rect 232222 50058 232306 50294
rect 232542 50058 232574 50294
rect 231954 14614 232574 50058
rect 231954 14378 231986 14614
rect 232222 14378 232306 14614
rect 232542 14378 232574 14614
rect 231954 14294 232574 14378
rect 231954 14058 231986 14294
rect 232222 14058 232306 14294
rect 232542 14058 232574 14294
rect 228234 -4422 228266 -4186
rect 228502 -4422 228586 -4186
rect 228822 -4422 228854 -4186
rect 228234 -4506 228854 -4422
rect 228234 -4742 228266 -4506
rect 228502 -4742 228586 -4506
rect 228822 -4742 228854 -4506
rect 228234 -5734 228854 -4742
rect 221954 -7302 221986 -7066
rect 222222 -7302 222306 -7066
rect 222542 -7302 222574 -7066
rect 221954 -7386 222574 -7302
rect 221954 -7622 221986 -7386
rect 222222 -7622 222306 -7386
rect 222542 -7622 222574 -7386
rect 221954 -7654 222574 -7622
rect 231954 -6106 232574 14058
rect 234514 707718 235134 707750
rect 234514 707482 234546 707718
rect 234782 707482 234866 707718
rect 235102 707482 235134 707718
rect 234514 707398 235134 707482
rect 234514 707162 234546 707398
rect 234782 707162 234866 707398
rect 235102 707162 235134 707398
rect 234514 673174 235134 707162
rect 234514 672938 234546 673174
rect 234782 672938 234866 673174
rect 235102 672938 235134 673174
rect 234514 672854 235134 672938
rect 234514 672618 234546 672854
rect 234782 672618 234866 672854
rect 235102 672618 235134 672854
rect 234514 637174 235134 672618
rect 234514 636938 234546 637174
rect 234782 636938 234866 637174
rect 235102 636938 235134 637174
rect 234514 636854 235134 636938
rect 234514 636618 234546 636854
rect 234782 636618 234866 636854
rect 235102 636618 235134 636854
rect 234514 601174 235134 636618
rect 234514 600938 234546 601174
rect 234782 600938 234866 601174
rect 235102 600938 235134 601174
rect 234514 600854 235134 600938
rect 234514 600618 234546 600854
rect 234782 600618 234866 600854
rect 235102 600618 235134 600854
rect 234514 565174 235134 600618
rect 234514 564938 234546 565174
rect 234782 564938 234866 565174
rect 235102 564938 235134 565174
rect 234514 564854 235134 564938
rect 234514 564618 234546 564854
rect 234782 564618 234866 564854
rect 235102 564618 235134 564854
rect 234514 529174 235134 564618
rect 234514 528938 234546 529174
rect 234782 528938 234866 529174
rect 235102 528938 235134 529174
rect 234514 528854 235134 528938
rect 234514 528618 234546 528854
rect 234782 528618 234866 528854
rect 235102 528618 235134 528854
rect 234514 493174 235134 528618
rect 234514 492938 234546 493174
rect 234782 492938 234866 493174
rect 235102 492938 235134 493174
rect 234514 492854 235134 492938
rect 234514 492618 234546 492854
rect 234782 492618 234866 492854
rect 235102 492618 235134 492854
rect 234514 457174 235134 492618
rect 234514 456938 234546 457174
rect 234782 456938 234866 457174
rect 235102 456938 235134 457174
rect 234514 456854 235134 456938
rect 234514 456618 234546 456854
rect 234782 456618 234866 456854
rect 235102 456618 235134 456854
rect 234514 421174 235134 456618
rect 234514 420938 234546 421174
rect 234782 420938 234866 421174
rect 235102 420938 235134 421174
rect 234514 420854 235134 420938
rect 234514 420618 234546 420854
rect 234782 420618 234866 420854
rect 235102 420618 235134 420854
rect 234514 385174 235134 420618
rect 234514 384938 234546 385174
rect 234782 384938 234866 385174
rect 235102 384938 235134 385174
rect 234514 384854 235134 384938
rect 234514 384618 234546 384854
rect 234782 384618 234866 384854
rect 235102 384618 235134 384854
rect 234514 349174 235134 384618
rect 234514 348938 234546 349174
rect 234782 348938 234866 349174
rect 235102 348938 235134 349174
rect 234514 348854 235134 348938
rect 234514 348618 234546 348854
rect 234782 348618 234866 348854
rect 235102 348618 235134 348854
rect 234514 313174 235134 348618
rect 234514 312938 234546 313174
rect 234782 312938 234866 313174
rect 235102 312938 235134 313174
rect 234514 312854 235134 312938
rect 234514 312618 234546 312854
rect 234782 312618 234866 312854
rect 235102 312618 235134 312854
rect 234514 277174 235134 312618
rect 234514 276938 234546 277174
rect 234782 276938 234866 277174
rect 235102 276938 235134 277174
rect 234514 276854 235134 276938
rect 234514 276618 234546 276854
rect 234782 276618 234866 276854
rect 235102 276618 235134 276854
rect 234514 241174 235134 276618
rect 234514 240938 234546 241174
rect 234782 240938 234866 241174
rect 235102 240938 235134 241174
rect 234514 240854 235134 240938
rect 234514 240618 234546 240854
rect 234782 240618 234866 240854
rect 235102 240618 235134 240854
rect 234514 205174 235134 240618
rect 234514 204938 234546 205174
rect 234782 204938 234866 205174
rect 235102 204938 235134 205174
rect 234514 204854 235134 204938
rect 234514 204618 234546 204854
rect 234782 204618 234866 204854
rect 235102 204618 235134 204854
rect 234514 169174 235134 204618
rect 234514 168938 234546 169174
rect 234782 168938 234866 169174
rect 235102 168938 235134 169174
rect 234514 168854 235134 168938
rect 234514 168618 234546 168854
rect 234782 168618 234866 168854
rect 235102 168618 235134 168854
rect 234514 133174 235134 168618
rect 234514 132938 234546 133174
rect 234782 132938 234866 133174
rect 235102 132938 235134 133174
rect 234514 132854 235134 132938
rect 234514 132618 234546 132854
rect 234782 132618 234866 132854
rect 235102 132618 235134 132854
rect 234514 97174 235134 132618
rect 234514 96938 234546 97174
rect 234782 96938 234866 97174
rect 235102 96938 235134 97174
rect 234514 96854 235134 96938
rect 234514 96618 234546 96854
rect 234782 96618 234866 96854
rect 235102 96618 235134 96854
rect 234514 61174 235134 96618
rect 234514 60938 234546 61174
rect 234782 60938 234866 61174
rect 235102 60938 235134 61174
rect 234514 60854 235134 60938
rect 234514 60618 234546 60854
rect 234782 60618 234866 60854
rect 235102 60618 235134 60854
rect 234514 25174 235134 60618
rect 234514 24938 234546 25174
rect 234782 24938 234866 25174
rect 235102 24938 235134 25174
rect 234514 24854 235134 24938
rect 234514 24618 234546 24854
rect 234782 24618 234866 24854
rect 235102 24618 235134 24854
rect 234514 -3226 235134 24618
rect 234514 -3462 234546 -3226
rect 234782 -3462 234866 -3226
rect 235102 -3462 235134 -3226
rect 234514 -3546 235134 -3462
rect 234514 -3782 234546 -3546
rect 234782 -3782 234866 -3546
rect 235102 -3782 235134 -3546
rect 234514 -3814 235134 -3782
rect 238234 676894 238854 709082
rect 238234 676658 238266 676894
rect 238502 676658 238586 676894
rect 238822 676658 238854 676894
rect 238234 676574 238854 676658
rect 238234 676338 238266 676574
rect 238502 676338 238586 676574
rect 238822 676338 238854 676574
rect 238234 640894 238854 676338
rect 238234 640658 238266 640894
rect 238502 640658 238586 640894
rect 238822 640658 238854 640894
rect 238234 640574 238854 640658
rect 238234 640338 238266 640574
rect 238502 640338 238586 640574
rect 238822 640338 238854 640574
rect 238234 604894 238854 640338
rect 238234 604658 238266 604894
rect 238502 604658 238586 604894
rect 238822 604658 238854 604894
rect 238234 604574 238854 604658
rect 238234 604338 238266 604574
rect 238502 604338 238586 604574
rect 238822 604338 238854 604574
rect 238234 568894 238854 604338
rect 238234 568658 238266 568894
rect 238502 568658 238586 568894
rect 238822 568658 238854 568894
rect 238234 568574 238854 568658
rect 238234 568338 238266 568574
rect 238502 568338 238586 568574
rect 238822 568338 238854 568574
rect 238234 532894 238854 568338
rect 238234 532658 238266 532894
rect 238502 532658 238586 532894
rect 238822 532658 238854 532894
rect 238234 532574 238854 532658
rect 238234 532338 238266 532574
rect 238502 532338 238586 532574
rect 238822 532338 238854 532574
rect 238234 496894 238854 532338
rect 238234 496658 238266 496894
rect 238502 496658 238586 496894
rect 238822 496658 238854 496894
rect 238234 496574 238854 496658
rect 238234 496338 238266 496574
rect 238502 496338 238586 496574
rect 238822 496338 238854 496574
rect 238234 460894 238854 496338
rect 238234 460658 238266 460894
rect 238502 460658 238586 460894
rect 238822 460658 238854 460894
rect 238234 460574 238854 460658
rect 238234 460338 238266 460574
rect 238502 460338 238586 460574
rect 238822 460338 238854 460574
rect 238234 424894 238854 460338
rect 238234 424658 238266 424894
rect 238502 424658 238586 424894
rect 238822 424658 238854 424894
rect 238234 424574 238854 424658
rect 238234 424338 238266 424574
rect 238502 424338 238586 424574
rect 238822 424338 238854 424574
rect 238234 388894 238854 424338
rect 238234 388658 238266 388894
rect 238502 388658 238586 388894
rect 238822 388658 238854 388894
rect 238234 388574 238854 388658
rect 238234 388338 238266 388574
rect 238502 388338 238586 388574
rect 238822 388338 238854 388574
rect 238234 352894 238854 388338
rect 238234 352658 238266 352894
rect 238502 352658 238586 352894
rect 238822 352658 238854 352894
rect 238234 352574 238854 352658
rect 238234 352338 238266 352574
rect 238502 352338 238586 352574
rect 238822 352338 238854 352574
rect 238234 316894 238854 352338
rect 238234 316658 238266 316894
rect 238502 316658 238586 316894
rect 238822 316658 238854 316894
rect 238234 316574 238854 316658
rect 238234 316338 238266 316574
rect 238502 316338 238586 316574
rect 238822 316338 238854 316574
rect 238234 280894 238854 316338
rect 238234 280658 238266 280894
rect 238502 280658 238586 280894
rect 238822 280658 238854 280894
rect 238234 280574 238854 280658
rect 238234 280338 238266 280574
rect 238502 280338 238586 280574
rect 238822 280338 238854 280574
rect 238234 244894 238854 280338
rect 238234 244658 238266 244894
rect 238502 244658 238586 244894
rect 238822 244658 238854 244894
rect 238234 244574 238854 244658
rect 238234 244338 238266 244574
rect 238502 244338 238586 244574
rect 238822 244338 238854 244574
rect 238234 208894 238854 244338
rect 238234 208658 238266 208894
rect 238502 208658 238586 208894
rect 238822 208658 238854 208894
rect 238234 208574 238854 208658
rect 238234 208338 238266 208574
rect 238502 208338 238586 208574
rect 238822 208338 238854 208574
rect 238234 172894 238854 208338
rect 238234 172658 238266 172894
rect 238502 172658 238586 172894
rect 238822 172658 238854 172894
rect 238234 172574 238854 172658
rect 238234 172338 238266 172574
rect 238502 172338 238586 172574
rect 238822 172338 238854 172574
rect 238234 136894 238854 172338
rect 238234 136658 238266 136894
rect 238502 136658 238586 136894
rect 238822 136658 238854 136894
rect 238234 136574 238854 136658
rect 238234 136338 238266 136574
rect 238502 136338 238586 136574
rect 238822 136338 238854 136574
rect 238234 100894 238854 136338
rect 238234 100658 238266 100894
rect 238502 100658 238586 100894
rect 238822 100658 238854 100894
rect 238234 100574 238854 100658
rect 238234 100338 238266 100574
rect 238502 100338 238586 100574
rect 238822 100338 238854 100574
rect 238234 64894 238854 100338
rect 238234 64658 238266 64894
rect 238502 64658 238586 64894
rect 238822 64658 238854 64894
rect 238234 64574 238854 64658
rect 238234 64338 238266 64574
rect 238502 64338 238586 64574
rect 238822 64338 238854 64574
rect 238234 28894 238854 64338
rect 238234 28658 238266 28894
rect 238502 28658 238586 28894
rect 238822 28658 238854 28894
rect 238234 28574 238854 28658
rect 238234 28338 238266 28574
rect 238502 28338 238586 28574
rect 238822 28338 238854 28574
rect 238234 -5146 238854 28338
rect 240794 704838 241414 705830
rect 240794 704602 240826 704838
rect 241062 704602 241146 704838
rect 241382 704602 241414 704838
rect 240794 704518 241414 704602
rect 240794 704282 240826 704518
rect 241062 704282 241146 704518
rect 241382 704282 241414 704518
rect 240794 687454 241414 704282
rect 240794 687218 240826 687454
rect 241062 687218 241146 687454
rect 241382 687218 241414 687454
rect 240794 687134 241414 687218
rect 240794 686898 240826 687134
rect 241062 686898 241146 687134
rect 241382 686898 241414 687134
rect 240794 651454 241414 686898
rect 240794 651218 240826 651454
rect 241062 651218 241146 651454
rect 241382 651218 241414 651454
rect 240794 651134 241414 651218
rect 240794 650898 240826 651134
rect 241062 650898 241146 651134
rect 241382 650898 241414 651134
rect 240794 615454 241414 650898
rect 240794 615218 240826 615454
rect 241062 615218 241146 615454
rect 241382 615218 241414 615454
rect 240794 615134 241414 615218
rect 240794 614898 240826 615134
rect 241062 614898 241146 615134
rect 241382 614898 241414 615134
rect 240794 579454 241414 614898
rect 240794 579218 240826 579454
rect 241062 579218 241146 579454
rect 241382 579218 241414 579454
rect 240794 579134 241414 579218
rect 240794 578898 240826 579134
rect 241062 578898 241146 579134
rect 241382 578898 241414 579134
rect 240794 543454 241414 578898
rect 240794 543218 240826 543454
rect 241062 543218 241146 543454
rect 241382 543218 241414 543454
rect 240794 543134 241414 543218
rect 240794 542898 240826 543134
rect 241062 542898 241146 543134
rect 241382 542898 241414 543134
rect 240794 507454 241414 542898
rect 240794 507218 240826 507454
rect 241062 507218 241146 507454
rect 241382 507218 241414 507454
rect 240794 507134 241414 507218
rect 240794 506898 240826 507134
rect 241062 506898 241146 507134
rect 241382 506898 241414 507134
rect 240794 471454 241414 506898
rect 240794 471218 240826 471454
rect 241062 471218 241146 471454
rect 241382 471218 241414 471454
rect 240794 471134 241414 471218
rect 240794 470898 240826 471134
rect 241062 470898 241146 471134
rect 241382 470898 241414 471134
rect 240794 435454 241414 470898
rect 240794 435218 240826 435454
rect 241062 435218 241146 435454
rect 241382 435218 241414 435454
rect 240794 435134 241414 435218
rect 240794 434898 240826 435134
rect 241062 434898 241146 435134
rect 241382 434898 241414 435134
rect 240794 399454 241414 434898
rect 240794 399218 240826 399454
rect 241062 399218 241146 399454
rect 241382 399218 241414 399454
rect 240794 399134 241414 399218
rect 240794 398898 240826 399134
rect 241062 398898 241146 399134
rect 241382 398898 241414 399134
rect 240794 363454 241414 398898
rect 240794 363218 240826 363454
rect 241062 363218 241146 363454
rect 241382 363218 241414 363454
rect 240794 363134 241414 363218
rect 240794 362898 240826 363134
rect 241062 362898 241146 363134
rect 241382 362898 241414 363134
rect 240794 327454 241414 362898
rect 240794 327218 240826 327454
rect 241062 327218 241146 327454
rect 241382 327218 241414 327454
rect 240794 327134 241414 327218
rect 240794 326898 240826 327134
rect 241062 326898 241146 327134
rect 241382 326898 241414 327134
rect 240794 291454 241414 326898
rect 240794 291218 240826 291454
rect 241062 291218 241146 291454
rect 241382 291218 241414 291454
rect 240794 291134 241414 291218
rect 240794 290898 240826 291134
rect 241062 290898 241146 291134
rect 241382 290898 241414 291134
rect 240794 255454 241414 290898
rect 240794 255218 240826 255454
rect 241062 255218 241146 255454
rect 241382 255218 241414 255454
rect 240794 255134 241414 255218
rect 240794 254898 240826 255134
rect 241062 254898 241146 255134
rect 241382 254898 241414 255134
rect 240794 219454 241414 254898
rect 240794 219218 240826 219454
rect 241062 219218 241146 219454
rect 241382 219218 241414 219454
rect 240794 219134 241414 219218
rect 240794 218898 240826 219134
rect 241062 218898 241146 219134
rect 241382 218898 241414 219134
rect 240794 183454 241414 218898
rect 240794 183218 240826 183454
rect 241062 183218 241146 183454
rect 241382 183218 241414 183454
rect 240794 183134 241414 183218
rect 240794 182898 240826 183134
rect 241062 182898 241146 183134
rect 241382 182898 241414 183134
rect 240794 147454 241414 182898
rect 240794 147218 240826 147454
rect 241062 147218 241146 147454
rect 241382 147218 241414 147454
rect 240794 147134 241414 147218
rect 240794 146898 240826 147134
rect 241062 146898 241146 147134
rect 241382 146898 241414 147134
rect 240794 111454 241414 146898
rect 240794 111218 240826 111454
rect 241062 111218 241146 111454
rect 241382 111218 241414 111454
rect 240794 111134 241414 111218
rect 240794 110898 240826 111134
rect 241062 110898 241146 111134
rect 241382 110898 241414 111134
rect 240794 75454 241414 110898
rect 240794 75218 240826 75454
rect 241062 75218 241146 75454
rect 241382 75218 241414 75454
rect 240794 75134 241414 75218
rect 240794 74898 240826 75134
rect 241062 74898 241146 75134
rect 241382 74898 241414 75134
rect 240794 39454 241414 74898
rect 240794 39218 240826 39454
rect 241062 39218 241146 39454
rect 241382 39218 241414 39454
rect 240794 39134 241414 39218
rect 240794 38898 240826 39134
rect 241062 38898 241146 39134
rect 241382 38898 241414 39134
rect 240794 3454 241414 38898
rect 240794 3218 240826 3454
rect 241062 3218 241146 3454
rect 241382 3218 241414 3454
rect 240794 3134 241414 3218
rect 240794 2898 240826 3134
rect 241062 2898 241146 3134
rect 241382 2898 241414 3134
rect 240794 -346 241414 2898
rect 240794 -582 240826 -346
rect 241062 -582 241146 -346
rect 241382 -582 241414 -346
rect 240794 -666 241414 -582
rect 240794 -902 240826 -666
rect 241062 -902 241146 -666
rect 241382 -902 241414 -666
rect 240794 -1894 241414 -902
rect 241954 680614 242574 711002
rect 251954 710598 252574 711590
rect 251954 710362 251986 710598
rect 252222 710362 252306 710598
rect 252542 710362 252574 710598
rect 251954 710278 252574 710362
rect 251954 710042 251986 710278
rect 252222 710042 252306 710278
rect 252542 710042 252574 710278
rect 248234 708678 248854 709670
rect 248234 708442 248266 708678
rect 248502 708442 248586 708678
rect 248822 708442 248854 708678
rect 248234 708358 248854 708442
rect 248234 708122 248266 708358
rect 248502 708122 248586 708358
rect 248822 708122 248854 708358
rect 241954 680378 241986 680614
rect 242222 680378 242306 680614
rect 242542 680378 242574 680614
rect 241954 680294 242574 680378
rect 241954 680058 241986 680294
rect 242222 680058 242306 680294
rect 242542 680058 242574 680294
rect 241954 644614 242574 680058
rect 241954 644378 241986 644614
rect 242222 644378 242306 644614
rect 242542 644378 242574 644614
rect 241954 644294 242574 644378
rect 241954 644058 241986 644294
rect 242222 644058 242306 644294
rect 242542 644058 242574 644294
rect 241954 608614 242574 644058
rect 241954 608378 241986 608614
rect 242222 608378 242306 608614
rect 242542 608378 242574 608614
rect 241954 608294 242574 608378
rect 241954 608058 241986 608294
rect 242222 608058 242306 608294
rect 242542 608058 242574 608294
rect 241954 572614 242574 608058
rect 241954 572378 241986 572614
rect 242222 572378 242306 572614
rect 242542 572378 242574 572614
rect 241954 572294 242574 572378
rect 241954 572058 241986 572294
rect 242222 572058 242306 572294
rect 242542 572058 242574 572294
rect 241954 536614 242574 572058
rect 241954 536378 241986 536614
rect 242222 536378 242306 536614
rect 242542 536378 242574 536614
rect 241954 536294 242574 536378
rect 241954 536058 241986 536294
rect 242222 536058 242306 536294
rect 242542 536058 242574 536294
rect 241954 500614 242574 536058
rect 241954 500378 241986 500614
rect 242222 500378 242306 500614
rect 242542 500378 242574 500614
rect 241954 500294 242574 500378
rect 241954 500058 241986 500294
rect 242222 500058 242306 500294
rect 242542 500058 242574 500294
rect 241954 464614 242574 500058
rect 241954 464378 241986 464614
rect 242222 464378 242306 464614
rect 242542 464378 242574 464614
rect 241954 464294 242574 464378
rect 241954 464058 241986 464294
rect 242222 464058 242306 464294
rect 242542 464058 242574 464294
rect 241954 428614 242574 464058
rect 241954 428378 241986 428614
rect 242222 428378 242306 428614
rect 242542 428378 242574 428614
rect 241954 428294 242574 428378
rect 241954 428058 241986 428294
rect 242222 428058 242306 428294
rect 242542 428058 242574 428294
rect 241954 392614 242574 428058
rect 241954 392378 241986 392614
rect 242222 392378 242306 392614
rect 242542 392378 242574 392614
rect 241954 392294 242574 392378
rect 241954 392058 241986 392294
rect 242222 392058 242306 392294
rect 242542 392058 242574 392294
rect 241954 356614 242574 392058
rect 241954 356378 241986 356614
rect 242222 356378 242306 356614
rect 242542 356378 242574 356614
rect 241954 356294 242574 356378
rect 241954 356058 241986 356294
rect 242222 356058 242306 356294
rect 242542 356058 242574 356294
rect 241954 320614 242574 356058
rect 241954 320378 241986 320614
rect 242222 320378 242306 320614
rect 242542 320378 242574 320614
rect 241954 320294 242574 320378
rect 241954 320058 241986 320294
rect 242222 320058 242306 320294
rect 242542 320058 242574 320294
rect 241954 284614 242574 320058
rect 241954 284378 241986 284614
rect 242222 284378 242306 284614
rect 242542 284378 242574 284614
rect 241954 284294 242574 284378
rect 241954 284058 241986 284294
rect 242222 284058 242306 284294
rect 242542 284058 242574 284294
rect 241954 248614 242574 284058
rect 241954 248378 241986 248614
rect 242222 248378 242306 248614
rect 242542 248378 242574 248614
rect 241954 248294 242574 248378
rect 241954 248058 241986 248294
rect 242222 248058 242306 248294
rect 242542 248058 242574 248294
rect 241954 212614 242574 248058
rect 241954 212378 241986 212614
rect 242222 212378 242306 212614
rect 242542 212378 242574 212614
rect 241954 212294 242574 212378
rect 241954 212058 241986 212294
rect 242222 212058 242306 212294
rect 242542 212058 242574 212294
rect 241954 176614 242574 212058
rect 241954 176378 241986 176614
rect 242222 176378 242306 176614
rect 242542 176378 242574 176614
rect 241954 176294 242574 176378
rect 241954 176058 241986 176294
rect 242222 176058 242306 176294
rect 242542 176058 242574 176294
rect 241954 140614 242574 176058
rect 241954 140378 241986 140614
rect 242222 140378 242306 140614
rect 242542 140378 242574 140614
rect 241954 140294 242574 140378
rect 241954 140058 241986 140294
rect 242222 140058 242306 140294
rect 242542 140058 242574 140294
rect 241954 104614 242574 140058
rect 241954 104378 241986 104614
rect 242222 104378 242306 104614
rect 242542 104378 242574 104614
rect 241954 104294 242574 104378
rect 241954 104058 241986 104294
rect 242222 104058 242306 104294
rect 242542 104058 242574 104294
rect 241954 68614 242574 104058
rect 241954 68378 241986 68614
rect 242222 68378 242306 68614
rect 242542 68378 242574 68614
rect 241954 68294 242574 68378
rect 241954 68058 241986 68294
rect 242222 68058 242306 68294
rect 242542 68058 242574 68294
rect 241954 32614 242574 68058
rect 241954 32378 241986 32614
rect 242222 32378 242306 32614
rect 242542 32378 242574 32614
rect 241954 32294 242574 32378
rect 241954 32058 241986 32294
rect 242222 32058 242306 32294
rect 242542 32058 242574 32294
rect 238234 -5382 238266 -5146
rect 238502 -5382 238586 -5146
rect 238822 -5382 238854 -5146
rect 238234 -5466 238854 -5382
rect 238234 -5702 238266 -5466
rect 238502 -5702 238586 -5466
rect 238822 -5702 238854 -5466
rect 238234 -5734 238854 -5702
rect 231954 -6342 231986 -6106
rect 232222 -6342 232306 -6106
rect 232542 -6342 232574 -6106
rect 231954 -6426 232574 -6342
rect 231954 -6662 231986 -6426
rect 232222 -6662 232306 -6426
rect 232542 -6662 232574 -6426
rect 231954 -7654 232574 -6662
rect 241954 -7066 242574 32058
rect 244514 706758 245134 707750
rect 244514 706522 244546 706758
rect 244782 706522 244866 706758
rect 245102 706522 245134 706758
rect 244514 706438 245134 706522
rect 244514 706202 244546 706438
rect 244782 706202 244866 706438
rect 245102 706202 245134 706438
rect 244514 691174 245134 706202
rect 244514 690938 244546 691174
rect 244782 690938 244866 691174
rect 245102 690938 245134 691174
rect 244514 690854 245134 690938
rect 244514 690618 244546 690854
rect 244782 690618 244866 690854
rect 245102 690618 245134 690854
rect 244514 655174 245134 690618
rect 244514 654938 244546 655174
rect 244782 654938 244866 655174
rect 245102 654938 245134 655174
rect 244514 654854 245134 654938
rect 244514 654618 244546 654854
rect 244782 654618 244866 654854
rect 245102 654618 245134 654854
rect 244514 619174 245134 654618
rect 244514 618938 244546 619174
rect 244782 618938 244866 619174
rect 245102 618938 245134 619174
rect 244514 618854 245134 618938
rect 244514 618618 244546 618854
rect 244782 618618 244866 618854
rect 245102 618618 245134 618854
rect 244514 583174 245134 618618
rect 244514 582938 244546 583174
rect 244782 582938 244866 583174
rect 245102 582938 245134 583174
rect 244514 582854 245134 582938
rect 244514 582618 244546 582854
rect 244782 582618 244866 582854
rect 245102 582618 245134 582854
rect 244514 547174 245134 582618
rect 244514 546938 244546 547174
rect 244782 546938 244866 547174
rect 245102 546938 245134 547174
rect 244514 546854 245134 546938
rect 244514 546618 244546 546854
rect 244782 546618 244866 546854
rect 245102 546618 245134 546854
rect 244514 511174 245134 546618
rect 244514 510938 244546 511174
rect 244782 510938 244866 511174
rect 245102 510938 245134 511174
rect 244514 510854 245134 510938
rect 244514 510618 244546 510854
rect 244782 510618 244866 510854
rect 245102 510618 245134 510854
rect 244514 475174 245134 510618
rect 244514 474938 244546 475174
rect 244782 474938 244866 475174
rect 245102 474938 245134 475174
rect 244514 474854 245134 474938
rect 244514 474618 244546 474854
rect 244782 474618 244866 474854
rect 245102 474618 245134 474854
rect 244514 439174 245134 474618
rect 244514 438938 244546 439174
rect 244782 438938 244866 439174
rect 245102 438938 245134 439174
rect 244514 438854 245134 438938
rect 244514 438618 244546 438854
rect 244782 438618 244866 438854
rect 245102 438618 245134 438854
rect 244514 403174 245134 438618
rect 244514 402938 244546 403174
rect 244782 402938 244866 403174
rect 245102 402938 245134 403174
rect 244514 402854 245134 402938
rect 244514 402618 244546 402854
rect 244782 402618 244866 402854
rect 245102 402618 245134 402854
rect 244514 367174 245134 402618
rect 244514 366938 244546 367174
rect 244782 366938 244866 367174
rect 245102 366938 245134 367174
rect 244514 366854 245134 366938
rect 244514 366618 244546 366854
rect 244782 366618 244866 366854
rect 245102 366618 245134 366854
rect 244514 331174 245134 366618
rect 244514 330938 244546 331174
rect 244782 330938 244866 331174
rect 245102 330938 245134 331174
rect 244514 330854 245134 330938
rect 244514 330618 244546 330854
rect 244782 330618 244866 330854
rect 245102 330618 245134 330854
rect 244514 295174 245134 330618
rect 244514 294938 244546 295174
rect 244782 294938 244866 295174
rect 245102 294938 245134 295174
rect 244514 294854 245134 294938
rect 244514 294618 244546 294854
rect 244782 294618 244866 294854
rect 245102 294618 245134 294854
rect 244514 259174 245134 294618
rect 244514 258938 244546 259174
rect 244782 258938 244866 259174
rect 245102 258938 245134 259174
rect 244514 258854 245134 258938
rect 244514 258618 244546 258854
rect 244782 258618 244866 258854
rect 245102 258618 245134 258854
rect 244514 223174 245134 258618
rect 244514 222938 244546 223174
rect 244782 222938 244866 223174
rect 245102 222938 245134 223174
rect 244514 222854 245134 222938
rect 244514 222618 244546 222854
rect 244782 222618 244866 222854
rect 245102 222618 245134 222854
rect 244514 187174 245134 222618
rect 244514 186938 244546 187174
rect 244782 186938 244866 187174
rect 245102 186938 245134 187174
rect 244514 186854 245134 186938
rect 244514 186618 244546 186854
rect 244782 186618 244866 186854
rect 245102 186618 245134 186854
rect 244514 151174 245134 186618
rect 244514 150938 244546 151174
rect 244782 150938 244866 151174
rect 245102 150938 245134 151174
rect 244514 150854 245134 150938
rect 244514 150618 244546 150854
rect 244782 150618 244866 150854
rect 245102 150618 245134 150854
rect 244514 115174 245134 150618
rect 244514 114938 244546 115174
rect 244782 114938 244866 115174
rect 245102 114938 245134 115174
rect 244514 114854 245134 114938
rect 244514 114618 244546 114854
rect 244782 114618 244866 114854
rect 245102 114618 245134 114854
rect 244514 79174 245134 114618
rect 244514 78938 244546 79174
rect 244782 78938 244866 79174
rect 245102 78938 245134 79174
rect 244514 78854 245134 78938
rect 244514 78618 244546 78854
rect 244782 78618 244866 78854
rect 245102 78618 245134 78854
rect 244514 43174 245134 78618
rect 244514 42938 244546 43174
rect 244782 42938 244866 43174
rect 245102 42938 245134 43174
rect 244514 42854 245134 42938
rect 244514 42618 244546 42854
rect 244782 42618 244866 42854
rect 245102 42618 245134 42854
rect 244514 7174 245134 42618
rect 244514 6938 244546 7174
rect 244782 6938 244866 7174
rect 245102 6938 245134 7174
rect 244514 6854 245134 6938
rect 244514 6618 244546 6854
rect 244782 6618 244866 6854
rect 245102 6618 245134 6854
rect 244514 -2266 245134 6618
rect 244514 -2502 244546 -2266
rect 244782 -2502 244866 -2266
rect 245102 -2502 245134 -2266
rect 244514 -2586 245134 -2502
rect 244514 -2822 244546 -2586
rect 244782 -2822 244866 -2586
rect 245102 -2822 245134 -2586
rect 244514 -3814 245134 -2822
rect 248234 694894 248854 708122
rect 248234 694658 248266 694894
rect 248502 694658 248586 694894
rect 248822 694658 248854 694894
rect 248234 694574 248854 694658
rect 248234 694338 248266 694574
rect 248502 694338 248586 694574
rect 248822 694338 248854 694574
rect 248234 658894 248854 694338
rect 248234 658658 248266 658894
rect 248502 658658 248586 658894
rect 248822 658658 248854 658894
rect 248234 658574 248854 658658
rect 248234 658338 248266 658574
rect 248502 658338 248586 658574
rect 248822 658338 248854 658574
rect 248234 622894 248854 658338
rect 248234 622658 248266 622894
rect 248502 622658 248586 622894
rect 248822 622658 248854 622894
rect 248234 622574 248854 622658
rect 248234 622338 248266 622574
rect 248502 622338 248586 622574
rect 248822 622338 248854 622574
rect 248234 586894 248854 622338
rect 248234 586658 248266 586894
rect 248502 586658 248586 586894
rect 248822 586658 248854 586894
rect 248234 586574 248854 586658
rect 248234 586338 248266 586574
rect 248502 586338 248586 586574
rect 248822 586338 248854 586574
rect 248234 550894 248854 586338
rect 248234 550658 248266 550894
rect 248502 550658 248586 550894
rect 248822 550658 248854 550894
rect 248234 550574 248854 550658
rect 248234 550338 248266 550574
rect 248502 550338 248586 550574
rect 248822 550338 248854 550574
rect 248234 514894 248854 550338
rect 248234 514658 248266 514894
rect 248502 514658 248586 514894
rect 248822 514658 248854 514894
rect 248234 514574 248854 514658
rect 248234 514338 248266 514574
rect 248502 514338 248586 514574
rect 248822 514338 248854 514574
rect 248234 478894 248854 514338
rect 248234 478658 248266 478894
rect 248502 478658 248586 478894
rect 248822 478658 248854 478894
rect 248234 478574 248854 478658
rect 248234 478338 248266 478574
rect 248502 478338 248586 478574
rect 248822 478338 248854 478574
rect 248234 442894 248854 478338
rect 248234 442658 248266 442894
rect 248502 442658 248586 442894
rect 248822 442658 248854 442894
rect 248234 442574 248854 442658
rect 248234 442338 248266 442574
rect 248502 442338 248586 442574
rect 248822 442338 248854 442574
rect 248234 406894 248854 442338
rect 248234 406658 248266 406894
rect 248502 406658 248586 406894
rect 248822 406658 248854 406894
rect 248234 406574 248854 406658
rect 248234 406338 248266 406574
rect 248502 406338 248586 406574
rect 248822 406338 248854 406574
rect 248234 370894 248854 406338
rect 248234 370658 248266 370894
rect 248502 370658 248586 370894
rect 248822 370658 248854 370894
rect 248234 370574 248854 370658
rect 248234 370338 248266 370574
rect 248502 370338 248586 370574
rect 248822 370338 248854 370574
rect 248234 334894 248854 370338
rect 248234 334658 248266 334894
rect 248502 334658 248586 334894
rect 248822 334658 248854 334894
rect 248234 334574 248854 334658
rect 248234 334338 248266 334574
rect 248502 334338 248586 334574
rect 248822 334338 248854 334574
rect 248234 298894 248854 334338
rect 248234 298658 248266 298894
rect 248502 298658 248586 298894
rect 248822 298658 248854 298894
rect 248234 298574 248854 298658
rect 248234 298338 248266 298574
rect 248502 298338 248586 298574
rect 248822 298338 248854 298574
rect 248234 262894 248854 298338
rect 248234 262658 248266 262894
rect 248502 262658 248586 262894
rect 248822 262658 248854 262894
rect 248234 262574 248854 262658
rect 248234 262338 248266 262574
rect 248502 262338 248586 262574
rect 248822 262338 248854 262574
rect 248234 226894 248854 262338
rect 248234 226658 248266 226894
rect 248502 226658 248586 226894
rect 248822 226658 248854 226894
rect 248234 226574 248854 226658
rect 248234 226338 248266 226574
rect 248502 226338 248586 226574
rect 248822 226338 248854 226574
rect 248234 190894 248854 226338
rect 248234 190658 248266 190894
rect 248502 190658 248586 190894
rect 248822 190658 248854 190894
rect 248234 190574 248854 190658
rect 248234 190338 248266 190574
rect 248502 190338 248586 190574
rect 248822 190338 248854 190574
rect 248234 154894 248854 190338
rect 248234 154658 248266 154894
rect 248502 154658 248586 154894
rect 248822 154658 248854 154894
rect 248234 154574 248854 154658
rect 248234 154338 248266 154574
rect 248502 154338 248586 154574
rect 248822 154338 248854 154574
rect 248234 118894 248854 154338
rect 248234 118658 248266 118894
rect 248502 118658 248586 118894
rect 248822 118658 248854 118894
rect 248234 118574 248854 118658
rect 248234 118338 248266 118574
rect 248502 118338 248586 118574
rect 248822 118338 248854 118574
rect 248234 82894 248854 118338
rect 248234 82658 248266 82894
rect 248502 82658 248586 82894
rect 248822 82658 248854 82894
rect 248234 82574 248854 82658
rect 248234 82338 248266 82574
rect 248502 82338 248586 82574
rect 248822 82338 248854 82574
rect 248234 46894 248854 82338
rect 248234 46658 248266 46894
rect 248502 46658 248586 46894
rect 248822 46658 248854 46894
rect 248234 46574 248854 46658
rect 248234 46338 248266 46574
rect 248502 46338 248586 46574
rect 248822 46338 248854 46574
rect 248234 10894 248854 46338
rect 248234 10658 248266 10894
rect 248502 10658 248586 10894
rect 248822 10658 248854 10894
rect 248234 10574 248854 10658
rect 248234 10338 248266 10574
rect 248502 10338 248586 10574
rect 248822 10338 248854 10574
rect 248234 -4186 248854 10338
rect 250794 705798 251414 705830
rect 250794 705562 250826 705798
rect 251062 705562 251146 705798
rect 251382 705562 251414 705798
rect 250794 705478 251414 705562
rect 250794 705242 250826 705478
rect 251062 705242 251146 705478
rect 251382 705242 251414 705478
rect 250794 669454 251414 705242
rect 250794 669218 250826 669454
rect 251062 669218 251146 669454
rect 251382 669218 251414 669454
rect 250794 669134 251414 669218
rect 250794 668898 250826 669134
rect 251062 668898 251146 669134
rect 251382 668898 251414 669134
rect 250794 633454 251414 668898
rect 250794 633218 250826 633454
rect 251062 633218 251146 633454
rect 251382 633218 251414 633454
rect 250794 633134 251414 633218
rect 250794 632898 250826 633134
rect 251062 632898 251146 633134
rect 251382 632898 251414 633134
rect 250794 597454 251414 632898
rect 250794 597218 250826 597454
rect 251062 597218 251146 597454
rect 251382 597218 251414 597454
rect 250794 597134 251414 597218
rect 250794 596898 250826 597134
rect 251062 596898 251146 597134
rect 251382 596898 251414 597134
rect 250794 561454 251414 596898
rect 250794 561218 250826 561454
rect 251062 561218 251146 561454
rect 251382 561218 251414 561454
rect 250794 561134 251414 561218
rect 250794 560898 250826 561134
rect 251062 560898 251146 561134
rect 251382 560898 251414 561134
rect 250794 525454 251414 560898
rect 250794 525218 250826 525454
rect 251062 525218 251146 525454
rect 251382 525218 251414 525454
rect 250794 525134 251414 525218
rect 250794 524898 250826 525134
rect 251062 524898 251146 525134
rect 251382 524898 251414 525134
rect 250794 489454 251414 524898
rect 250794 489218 250826 489454
rect 251062 489218 251146 489454
rect 251382 489218 251414 489454
rect 250794 489134 251414 489218
rect 250794 488898 250826 489134
rect 251062 488898 251146 489134
rect 251382 488898 251414 489134
rect 250794 453454 251414 488898
rect 250794 453218 250826 453454
rect 251062 453218 251146 453454
rect 251382 453218 251414 453454
rect 250794 453134 251414 453218
rect 250794 452898 250826 453134
rect 251062 452898 251146 453134
rect 251382 452898 251414 453134
rect 250794 417454 251414 452898
rect 250794 417218 250826 417454
rect 251062 417218 251146 417454
rect 251382 417218 251414 417454
rect 250794 417134 251414 417218
rect 250794 416898 250826 417134
rect 251062 416898 251146 417134
rect 251382 416898 251414 417134
rect 250794 381454 251414 416898
rect 250794 381218 250826 381454
rect 251062 381218 251146 381454
rect 251382 381218 251414 381454
rect 250794 381134 251414 381218
rect 250794 380898 250826 381134
rect 251062 380898 251146 381134
rect 251382 380898 251414 381134
rect 250794 345454 251414 380898
rect 250794 345218 250826 345454
rect 251062 345218 251146 345454
rect 251382 345218 251414 345454
rect 250794 345134 251414 345218
rect 250794 344898 250826 345134
rect 251062 344898 251146 345134
rect 251382 344898 251414 345134
rect 250794 309454 251414 344898
rect 250794 309218 250826 309454
rect 251062 309218 251146 309454
rect 251382 309218 251414 309454
rect 250794 309134 251414 309218
rect 250794 308898 250826 309134
rect 251062 308898 251146 309134
rect 251382 308898 251414 309134
rect 250794 273454 251414 308898
rect 250794 273218 250826 273454
rect 251062 273218 251146 273454
rect 251382 273218 251414 273454
rect 250794 273134 251414 273218
rect 250794 272898 250826 273134
rect 251062 272898 251146 273134
rect 251382 272898 251414 273134
rect 250794 237454 251414 272898
rect 250794 237218 250826 237454
rect 251062 237218 251146 237454
rect 251382 237218 251414 237454
rect 250794 237134 251414 237218
rect 250794 236898 250826 237134
rect 251062 236898 251146 237134
rect 251382 236898 251414 237134
rect 250794 201454 251414 236898
rect 250794 201218 250826 201454
rect 251062 201218 251146 201454
rect 251382 201218 251414 201454
rect 250794 201134 251414 201218
rect 250794 200898 250826 201134
rect 251062 200898 251146 201134
rect 251382 200898 251414 201134
rect 250794 165454 251414 200898
rect 250794 165218 250826 165454
rect 251062 165218 251146 165454
rect 251382 165218 251414 165454
rect 250794 165134 251414 165218
rect 250794 164898 250826 165134
rect 251062 164898 251146 165134
rect 251382 164898 251414 165134
rect 250794 129454 251414 164898
rect 250794 129218 250826 129454
rect 251062 129218 251146 129454
rect 251382 129218 251414 129454
rect 250794 129134 251414 129218
rect 250794 128898 250826 129134
rect 251062 128898 251146 129134
rect 251382 128898 251414 129134
rect 250794 93454 251414 128898
rect 250794 93218 250826 93454
rect 251062 93218 251146 93454
rect 251382 93218 251414 93454
rect 250794 93134 251414 93218
rect 250794 92898 250826 93134
rect 251062 92898 251146 93134
rect 251382 92898 251414 93134
rect 250794 57454 251414 92898
rect 250794 57218 250826 57454
rect 251062 57218 251146 57454
rect 251382 57218 251414 57454
rect 250794 57134 251414 57218
rect 250794 56898 250826 57134
rect 251062 56898 251146 57134
rect 251382 56898 251414 57134
rect 250794 21454 251414 56898
rect 250794 21218 250826 21454
rect 251062 21218 251146 21454
rect 251382 21218 251414 21454
rect 250794 21134 251414 21218
rect 250794 20898 250826 21134
rect 251062 20898 251146 21134
rect 251382 20898 251414 21134
rect 250794 -1306 251414 20898
rect 250794 -1542 250826 -1306
rect 251062 -1542 251146 -1306
rect 251382 -1542 251414 -1306
rect 250794 -1626 251414 -1542
rect 250794 -1862 250826 -1626
rect 251062 -1862 251146 -1626
rect 251382 -1862 251414 -1626
rect 250794 -1894 251414 -1862
rect 251954 698614 252574 710042
rect 261954 711558 262574 711590
rect 261954 711322 261986 711558
rect 262222 711322 262306 711558
rect 262542 711322 262574 711558
rect 261954 711238 262574 711322
rect 261954 711002 261986 711238
rect 262222 711002 262306 711238
rect 262542 711002 262574 711238
rect 258234 709638 258854 709670
rect 258234 709402 258266 709638
rect 258502 709402 258586 709638
rect 258822 709402 258854 709638
rect 258234 709318 258854 709402
rect 258234 709082 258266 709318
rect 258502 709082 258586 709318
rect 258822 709082 258854 709318
rect 251954 698378 251986 698614
rect 252222 698378 252306 698614
rect 252542 698378 252574 698614
rect 251954 698294 252574 698378
rect 251954 698058 251986 698294
rect 252222 698058 252306 698294
rect 252542 698058 252574 698294
rect 251954 662614 252574 698058
rect 251954 662378 251986 662614
rect 252222 662378 252306 662614
rect 252542 662378 252574 662614
rect 251954 662294 252574 662378
rect 251954 662058 251986 662294
rect 252222 662058 252306 662294
rect 252542 662058 252574 662294
rect 251954 626614 252574 662058
rect 251954 626378 251986 626614
rect 252222 626378 252306 626614
rect 252542 626378 252574 626614
rect 251954 626294 252574 626378
rect 251954 626058 251986 626294
rect 252222 626058 252306 626294
rect 252542 626058 252574 626294
rect 251954 590614 252574 626058
rect 251954 590378 251986 590614
rect 252222 590378 252306 590614
rect 252542 590378 252574 590614
rect 251954 590294 252574 590378
rect 251954 590058 251986 590294
rect 252222 590058 252306 590294
rect 252542 590058 252574 590294
rect 251954 554614 252574 590058
rect 251954 554378 251986 554614
rect 252222 554378 252306 554614
rect 252542 554378 252574 554614
rect 251954 554294 252574 554378
rect 251954 554058 251986 554294
rect 252222 554058 252306 554294
rect 252542 554058 252574 554294
rect 251954 518614 252574 554058
rect 251954 518378 251986 518614
rect 252222 518378 252306 518614
rect 252542 518378 252574 518614
rect 251954 518294 252574 518378
rect 251954 518058 251986 518294
rect 252222 518058 252306 518294
rect 252542 518058 252574 518294
rect 251954 482614 252574 518058
rect 251954 482378 251986 482614
rect 252222 482378 252306 482614
rect 252542 482378 252574 482614
rect 251954 482294 252574 482378
rect 251954 482058 251986 482294
rect 252222 482058 252306 482294
rect 252542 482058 252574 482294
rect 251954 446614 252574 482058
rect 251954 446378 251986 446614
rect 252222 446378 252306 446614
rect 252542 446378 252574 446614
rect 251954 446294 252574 446378
rect 251954 446058 251986 446294
rect 252222 446058 252306 446294
rect 252542 446058 252574 446294
rect 251954 410614 252574 446058
rect 251954 410378 251986 410614
rect 252222 410378 252306 410614
rect 252542 410378 252574 410614
rect 251954 410294 252574 410378
rect 251954 410058 251986 410294
rect 252222 410058 252306 410294
rect 252542 410058 252574 410294
rect 251954 374614 252574 410058
rect 251954 374378 251986 374614
rect 252222 374378 252306 374614
rect 252542 374378 252574 374614
rect 251954 374294 252574 374378
rect 251954 374058 251986 374294
rect 252222 374058 252306 374294
rect 252542 374058 252574 374294
rect 251954 338614 252574 374058
rect 251954 338378 251986 338614
rect 252222 338378 252306 338614
rect 252542 338378 252574 338614
rect 251954 338294 252574 338378
rect 251954 338058 251986 338294
rect 252222 338058 252306 338294
rect 252542 338058 252574 338294
rect 251954 302614 252574 338058
rect 251954 302378 251986 302614
rect 252222 302378 252306 302614
rect 252542 302378 252574 302614
rect 251954 302294 252574 302378
rect 251954 302058 251986 302294
rect 252222 302058 252306 302294
rect 252542 302058 252574 302294
rect 251954 266614 252574 302058
rect 251954 266378 251986 266614
rect 252222 266378 252306 266614
rect 252542 266378 252574 266614
rect 251954 266294 252574 266378
rect 251954 266058 251986 266294
rect 252222 266058 252306 266294
rect 252542 266058 252574 266294
rect 251954 230614 252574 266058
rect 251954 230378 251986 230614
rect 252222 230378 252306 230614
rect 252542 230378 252574 230614
rect 251954 230294 252574 230378
rect 251954 230058 251986 230294
rect 252222 230058 252306 230294
rect 252542 230058 252574 230294
rect 251954 194614 252574 230058
rect 251954 194378 251986 194614
rect 252222 194378 252306 194614
rect 252542 194378 252574 194614
rect 251954 194294 252574 194378
rect 251954 194058 251986 194294
rect 252222 194058 252306 194294
rect 252542 194058 252574 194294
rect 251954 158614 252574 194058
rect 251954 158378 251986 158614
rect 252222 158378 252306 158614
rect 252542 158378 252574 158614
rect 251954 158294 252574 158378
rect 251954 158058 251986 158294
rect 252222 158058 252306 158294
rect 252542 158058 252574 158294
rect 251954 122614 252574 158058
rect 251954 122378 251986 122614
rect 252222 122378 252306 122614
rect 252542 122378 252574 122614
rect 251954 122294 252574 122378
rect 251954 122058 251986 122294
rect 252222 122058 252306 122294
rect 252542 122058 252574 122294
rect 251954 86614 252574 122058
rect 251954 86378 251986 86614
rect 252222 86378 252306 86614
rect 252542 86378 252574 86614
rect 251954 86294 252574 86378
rect 251954 86058 251986 86294
rect 252222 86058 252306 86294
rect 252542 86058 252574 86294
rect 251954 50614 252574 86058
rect 251954 50378 251986 50614
rect 252222 50378 252306 50614
rect 252542 50378 252574 50614
rect 251954 50294 252574 50378
rect 251954 50058 251986 50294
rect 252222 50058 252306 50294
rect 252542 50058 252574 50294
rect 251954 14614 252574 50058
rect 251954 14378 251986 14614
rect 252222 14378 252306 14614
rect 252542 14378 252574 14614
rect 251954 14294 252574 14378
rect 251954 14058 251986 14294
rect 252222 14058 252306 14294
rect 252542 14058 252574 14294
rect 248234 -4422 248266 -4186
rect 248502 -4422 248586 -4186
rect 248822 -4422 248854 -4186
rect 248234 -4506 248854 -4422
rect 248234 -4742 248266 -4506
rect 248502 -4742 248586 -4506
rect 248822 -4742 248854 -4506
rect 248234 -5734 248854 -4742
rect 241954 -7302 241986 -7066
rect 242222 -7302 242306 -7066
rect 242542 -7302 242574 -7066
rect 241954 -7386 242574 -7302
rect 241954 -7622 241986 -7386
rect 242222 -7622 242306 -7386
rect 242542 -7622 242574 -7386
rect 241954 -7654 242574 -7622
rect 251954 -6106 252574 14058
rect 254514 707718 255134 707750
rect 254514 707482 254546 707718
rect 254782 707482 254866 707718
rect 255102 707482 255134 707718
rect 254514 707398 255134 707482
rect 254514 707162 254546 707398
rect 254782 707162 254866 707398
rect 255102 707162 255134 707398
rect 254514 673174 255134 707162
rect 254514 672938 254546 673174
rect 254782 672938 254866 673174
rect 255102 672938 255134 673174
rect 254514 672854 255134 672938
rect 254514 672618 254546 672854
rect 254782 672618 254866 672854
rect 255102 672618 255134 672854
rect 254514 637174 255134 672618
rect 254514 636938 254546 637174
rect 254782 636938 254866 637174
rect 255102 636938 255134 637174
rect 254514 636854 255134 636938
rect 254514 636618 254546 636854
rect 254782 636618 254866 636854
rect 255102 636618 255134 636854
rect 254514 601174 255134 636618
rect 254514 600938 254546 601174
rect 254782 600938 254866 601174
rect 255102 600938 255134 601174
rect 254514 600854 255134 600938
rect 254514 600618 254546 600854
rect 254782 600618 254866 600854
rect 255102 600618 255134 600854
rect 254514 565174 255134 600618
rect 254514 564938 254546 565174
rect 254782 564938 254866 565174
rect 255102 564938 255134 565174
rect 254514 564854 255134 564938
rect 254514 564618 254546 564854
rect 254782 564618 254866 564854
rect 255102 564618 255134 564854
rect 254514 529174 255134 564618
rect 254514 528938 254546 529174
rect 254782 528938 254866 529174
rect 255102 528938 255134 529174
rect 254514 528854 255134 528938
rect 254514 528618 254546 528854
rect 254782 528618 254866 528854
rect 255102 528618 255134 528854
rect 254514 493174 255134 528618
rect 254514 492938 254546 493174
rect 254782 492938 254866 493174
rect 255102 492938 255134 493174
rect 254514 492854 255134 492938
rect 254514 492618 254546 492854
rect 254782 492618 254866 492854
rect 255102 492618 255134 492854
rect 254514 457174 255134 492618
rect 254514 456938 254546 457174
rect 254782 456938 254866 457174
rect 255102 456938 255134 457174
rect 254514 456854 255134 456938
rect 254514 456618 254546 456854
rect 254782 456618 254866 456854
rect 255102 456618 255134 456854
rect 254514 421174 255134 456618
rect 254514 420938 254546 421174
rect 254782 420938 254866 421174
rect 255102 420938 255134 421174
rect 254514 420854 255134 420938
rect 254514 420618 254546 420854
rect 254782 420618 254866 420854
rect 255102 420618 255134 420854
rect 254514 385174 255134 420618
rect 254514 384938 254546 385174
rect 254782 384938 254866 385174
rect 255102 384938 255134 385174
rect 254514 384854 255134 384938
rect 254514 384618 254546 384854
rect 254782 384618 254866 384854
rect 255102 384618 255134 384854
rect 254514 349174 255134 384618
rect 254514 348938 254546 349174
rect 254782 348938 254866 349174
rect 255102 348938 255134 349174
rect 254514 348854 255134 348938
rect 254514 348618 254546 348854
rect 254782 348618 254866 348854
rect 255102 348618 255134 348854
rect 254514 313174 255134 348618
rect 254514 312938 254546 313174
rect 254782 312938 254866 313174
rect 255102 312938 255134 313174
rect 254514 312854 255134 312938
rect 254514 312618 254546 312854
rect 254782 312618 254866 312854
rect 255102 312618 255134 312854
rect 254514 277174 255134 312618
rect 254514 276938 254546 277174
rect 254782 276938 254866 277174
rect 255102 276938 255134 277174
rect 254514 276854 255134 276938
rect 254514 276618 254546 276854
rect 254782 276618 254866 276854
rect 255102 276618 255134 276854
rect 254514 241174 255134 276618
rect 254514 240938 254546 241174
rect 254782 240938 254866 241174
rect 255102 240938 255134 241174
rect 254514 240854 255134 240938
rect 254514 240618 254546 240854
rect 254782 240618 254866 240854
rect 255102 240618 255134 240854
rect 254514 205174 255134 240618
rect 254514 204938 254546 205174
rect 254782 204938 254866 205174
rect 255102 204938 255134 205174
rect 254514 204854 255134 204938
rect 254514 204618 254546 204854
rect 254782 204618 254866 204854
rect 255102 204618 255134 204854
rect 254514 169174 255134 204618
rect 254514 168938 254546 169174
rect 254782 168938 254866 169174
rect 255102 168938 255134 169174
rect 254514 168854 255134 168938
rect 254514 168618 254546 168854
rect 254782 168618 254866 168854
rect 255102 168618 255134 168854
rect 254514 133174 255134 168618
rect 254514 132938 254546 133174
rect 254782 132938 254866 133174
rect 255102 132938 255134 133174
rect 254514 132854 255134 132938
rect 254514 132618 254546 132854
rect 254782 132618 254866 132854
rect 255102 132618 255134 132854
rect 254514 97174 255134 132618
rect 254514 96938 254546 97174
rect 254782 96938 254866 97174
rect 255102 96938 255134 97174
rect 254514 96854 255134 96938
rect 254514 96618 254546 96854
rect 254782 96618 254866 96854
rect 255102 96618 255134 96854
rect 254514 61174 255134 96618
rect 254514 60938 254546 61174
rect 254782 60938 254866 61174
rect 255102 60938 255134 61174
rect 254514 60854 255134 60938
rect 254514 60618 254546 60854
rect 254782 60618 254866 60854
rect 255102 60618 255134 60854
rect 254514 25174 255134 60618
rect 254514 24938 254546 25174
rect 254782 24938 254866 25174
rect 255102 24938 255134 25174
rect 254514 24854 255134 24938
rect 254514 24618 254546 24854
rect 254782 24618 254866 24854
rect 255102 24618 255134 24854
rect 254514 -3226 255134 24618
rect 254514 -3462 254546 -3226
rect 254782 -3462 254866 -3226
rect 255102 -3462 255134 -3226
rect 254514 -3546 255134 -3462
rect 254514 -3782 254546 -3546
rect 254782 -3782 254866 -3546
rect 255102 -3782 255134 -3546
rect 254514 -3814 255134 -3782
rect 258234 676894 258854 709082
rect 258234 676658 258266 676894
rect 258502 676658 258586 676894
rect 258822 676658 258854 676894
rect 258234 676574 258854 676658
rect 258234 676338 258266 676574
rect 258502 676338 258586 676574
rect 258822 676338 258854 676574
rect 258234 640894 258854 676338
rect 258234 640658 258266 640894
rect 258502 640658 258586 640894
rect 258822 640658 258854 640894
rect 258234 640574 258854 640658
rect 258234 640338 258266 640574
rect 258502 640338 258586 640574
rect 258822 640338 258854 640574
rect 258234 604894 258854 640338
rect 258234 604658 258266 604894
rect 258502 604658 258586 604894
rect 258822 604658 258854 604894
rect 258234 604574 258854 604658
rect 258234 604338 258266 604574
rect 258502 604338 258586 604574
rect 258822 604338 258854 604574
rect 258234 568894 258854 604338
rect 258234 568658 258266 568894
rect 258502 568658 258586 568894
rect 258822 568658 258854 568894
rect 258234 568574 258854 568658
rect 258234 568338 258266 568574
rect 258502 568338 258586 568574
rect 258822 568338 258854 568574
rect 258234 532894 258854 568338
rect 258234 532658 258266 532894
rect 258502 532658 258586 532894
rect 258822 532658 258854 532894
rect 258234 532574 258854 532658
rect 258234 532338 258266 532574
rect 258502 532338 258586 532574
rect 258822 532338 258854 532574
rect 258234 496894 258854 532338
rect 258234 496658 258266 496894
rect 258502 496658 258586 496894
rect 258822 496658 258854 496894
rect 258234 496574 258854 496658
rect 258234 496338 258266 496574
rect 258502 496338 258586 496574
rect 258822 496338 258854 496574
rect 258234 460894 258854 496338
rect 258234 460658 258266 460894
rect 258502 460658 258586 460894
rect 258822 460658 258854 460894
rect 258234 460574 258854 460658
rect 258234 460338 258266 460574
rect 258502 460338 258586 460574
rect 258822 460338 258854 460574
rect 258234 424894 258854 460338
rect 258234 424658 258266 424894
rect 258502 424658 258586 424894
rect 258822 424658 258854 424894
rect 258234 424574 258854 424658
rect 258234 424338 258266 424574
rect 258502 424338 258586 424574
rect 258822 424338 258854 424574
rect 258234 388894 258854 424338
rect 258234 388658 258266 388894
rect 258502 388658 258586 388894
rect 258822 388658 258854 388894
rect 258234 388574 258854 388658
rect 258234 388338 258266 388574
rect 258502 388338 258586 388574
rect 258822 388338 258854 388574
rect 258234 352894 258854 388338
rect 258234 352658 258266 352894
rect 258502 352658 258586 352894
rect 258822 352658 258854 352894
rect 258234 352574 258854 352658
rect 258234 352338 258266 352574
rect 258502 352338 258586 352574
rect 258822 352338 258854 352574
rect 258234 316894 258854 352338
rect 258234 316658 258266 316894
rect 258502 316658 258586 316894
rect 258822 316658 258854 316894
rect 258234 316574 258854 316658
rect 258234 316338 258266 316574
rect 258502 316338 258586 316574
rect 258822 316338 258854 316574
rect 258234 280894 258854 316338
rect 258234 280658 258266 280894
rect 258502 280658 258586 280894
rect 258822 280658 258854 280894
rect 258234 280574 258854 280658
rect 258234 280338 258266 280574
rect 258502 280338 258586 280574
rect 258822 280338 258854 280574
rect 258234 244894 258854 280338
rect 258234 244658 258266 244894
rect 258502 244658 258586 244894
rect 258822 244658 258854 244894
rect 258234 244574 258854 244658
rect 258234 244338 258266 244574
rect 258502 244338 258586 244574
rect 258822 244338 258854 244574
rect 258234 208894 258854 244338
rect 258234 208658 258266 208894
rect 258502 208658 258586 208894
rect 258822 208658 258854 208894
rect 258234 208574 258854 208658
rect 258234 208338 258266 208574
rect 258502 208338 258586 208574
rect 258822 208338 258854 208574
rect 258234 172894 258854 208338
rect 258234 172658 258266 172894
rect 258502 172658 258586 172894
rect 258822 172658 258854 172894
rect 258234 172574 258854 172658
rect 258234 172338 258266 172574
rect 258502 172338 258586 172574
rect 258822 172338 258854 172574
rect 258234 136894 258854 172338
rect 258234 136658 258266 136894
rect 258502 136658 258586 136894
rect 258822 136658 258854 136894
rect 258234 136574 258854 136658
rect 258234 136338 258266 136574
rect 258502 136338 258586 136574
rect 258822 136338 258854 136574
rect 258234 100894 258854 136338
rect 258234 100658 258266 100894
rect 258502 100658 258586 100894
rect 258822 100658 258854 100894
rect 258234 100574 258854 100658
rect 258234 100338 258266 100574
rect 258502 100338 258586 100574
rect 258822 100338 258854 100574
rect 258234 64894 258854 100338
rect 258234 64658 258266 64894
rect 258502 64658 258586 64894
rect 258822 64658 258854 64894
rect 258234 64574 258854 64658
rect 258234 64338 258266 64574
rect 258502 64338 258586 64574
rect 258822 64338 258854 64574
rect 258234 28894 258854 64338
rect 258234 28658 258266 28894
rect 258502 28658 258586 28894
rect 258822 28658 258854 28894
rect 258234 28574 258854 28658
rect 258234 28338 258266 28574
rect 258502 28338 258586 28574
rect 258822 28338 258854 28574
rect 258234 -5146 258854 28338
rect 260794 704838 261414 705830
rect 260794 704602 260826 704838
rect 261062 704602 261146 704838
rect 261382 704602 261414 704838
rect 260794 704518 261414 704602
rect 260794 704282 260826 704518
rect 261062 704282 261146 704518
rect 261382 704282 261414 704518
rect 260794 687454 261414 704282
rect 260794 687218 260826 687454
rect 261062 687218 261146 687454
rect 261382 687218 261414 687454
rect 260794 687134 261414 687218
rect 260794 686898 260826 687134
rect 261062 686898 261146 687134
rect 261382 686898 261414 687134
rect 260794 651454 261414 686898
rect 260794 651218 260826 651454
rect 261062 651218 261146 651454
rect 261382 651218 261414 651454
rect 260794 651134 261414 651218
rect 260794 650898 260826 651134
rect 261062 650898 261146 651134
rect 261382 650898 261414 651134
rect 260794 615454 261414 650898
rect 260794 615218 260826 615454
rect 261062 615218 261146 615454
rect 261382 615218 261414 615454
rect 260794 615134 261414 615218
rect 260794 614898 260826 615134
rect 261062 614898 261146 615134
rect 261382 614898 261414 615134
rect 260794 579454 261414 614898
rect 260794 579218 260826 579454
rect 261062 579218 261146 579454
rect 261382 579218 261414 579454
rect 260794 579134 261414 579218
rect 260794 578898 260826 579134
rect 261062 578898 261146 579134
rect 261382 578898 261414 579134
rect 260794 543454 261414 578898
rect 260794 543218 260826 543454
rect 261062 543218 261146 543454
rect 261382 543218 261414 543454
rect 260794 543134 261414 543218
rect 260794 542898 260826 543134
rect 261062 542898 261146 543134
rect 261382 542898 261414 543134
rect 260794 507454 261414 542898
rect 260794 507218 260826 507454
rect 261062 507218 261146 507454
rect 261382 507218 261414 507454
rect 260794 507134 261414 507218
rect 260794 506898 260826 507134
rect 261062 506898 261146 507134
rect 261382 506898 261414 507134
rect 260794 471454 261414 506898
rect 260794 471218 260826 471454
rect 261062 471218 261146 471454
rect 261382 471218 261414 471454
rect 260794 471134 261414 471218
rect 260794 470898 260826 471134
rect 261062 470898 261146 471134
rect 261382 470898 261414 471134
rect 260794 435454 261414 470898
rect 260794 435218 260826 435454
rect 261062 435218 261146 435454
rect 261382 435218 261414 435454
rect 260794 435134 261414 435218
rect 260794 434898 260826 435134
rect 261062 434898 261146 435134
rect 261382 434898 261414 435134
rect 260794 399454 261414 434898
rect 260794 399218 260826 399454
rect 261062 399218 261146 399454
rect 261382 399218 261414 399454
rect 260794 399134 261414 399218
rect 260794 398898 260826 399134
rect 261062 398898 261146 399134
rect 261382 398898 261414 399134
rect 260794 363454 261414 398898
rect 260794 363218 260826 363454
rect 261062 363218 261146 363454
rect 261382 363218 261414 363454
rect 260794 363134 261414 363218
rect 260794 362898 260826 363134
rect 261062 362898 261146 363134
rect 261382 362898 261414 363134
rect 260794 327454 261414 362898
rect 260794 327218 260826 327454
rect 261062 327218 261146 327454
rect 261382 327218 261414 327454
rect 260794 327134 261414 327218
rect 260794 326898 260826 327134
rect 261062 326898 261146 327134
rect 261382 326898 261414 327134
rect 260794 291454 261414 326898
rect 260794 291218 260826 291454
rect 261062 291218 261146 291454
rect 261382 291218 261414 291454
rect 260794 291134 261414 291218
rect 260794 290898 260826 291134
rect 261062 290898 261146 291134
rect 261382 290898 261414 291134
rect 260794 255454 261414 290898
rect 260794 255218 260826 255454
rect 261062 255218 261146 255454
rect 261382 255218 261414 255454
rect 260794 255134 261414 255218
rect 260794 254898 260826 255134
rect 261062 254898 261146 255134
rect 261382 254898 261414 255134
rect 260794 219454 261414 254898
rect 260794 219218 260826 219454
rect 261062 219218 261146 219454
rect 261382 219218 261414 219454
rect 260794 219134 261414 219218
rect 260794 218898 260826 219134
rect 261062 218898 261146 219134
rect 261382 218898 261414 219134
rect 260794 183454 261414 218898
rect 260794 183218 260826 183454
rect 261062 183218 261146 183454
rect 261382 183218 261414 183454
rect 260794 183134 261414 183218
rect 260794 182898 260826 183134
rect 261062 182898 261146 183134
rect 261382 182898 261414 183134
rect 260794 147454 261414 182898
rect 260794 147218 260826 147454
rect 261062 147218 261146 147454
rect 261382 147218 261414 147454
rect 260794 147134 261414 147218
rect 260794 146898 260826 147134
rect 261062 146898 261146 147134
rect 261382 146898 261414 147134
rect 260794 111454 261414 146898
rect 260794 111218 260826 111454
rect 261062 111218 261146 111454
rect 261382 111218 261414 111454
rect 260794 111134 261414 111218
rect 260794 110898 260826 111134
rect 261062 110898 261146 111134
rect 261382 110898 261414 111134
rect 260794 75454 261414 110898
rect 260794 75218 260826 75454
rect 261062 75218 261146 75454
rect 261382 75218 261414 75454
rect 260794 75134 261414 75218
rect 260794 74898 260826 75134
rect 261062 74898 261146 75134
rect 261382 74898 261414 75134
rect 260794 39454 261414 74898
rect 260794 39218 260826 39454
rect 261062 39218 261146 39454
rect 261382 39218 261414 39454
rect 260794 39134 261414 39218
rect 260794 38898 260826 39134
rect 261062 38898 261146 39134
rect 261382 38898 261414 39134
rect 260794 3454 261414 38898
rect 260794 3218 260826 3454
rect 261062 3218 261146 3454
rect 261382 3218 261414 3454
rect 260794 3134 261414 3218
rect 260794 2898 260826 3134
rect 261062 2898 261146 3134
rect 261382 2898 261414 3134
rect 260794 -346 261414 2898
rect 260794 -582 260826 -346
rect 261062 -582 261146 -346
rect 261382 -582 261414 -346
rect 260794 -666 261414 -582
rect 260794 -902 260826 -666
rect 261062 -902 261146 -666
rect 261382 -902 261414 -666
rect 260794 -1894 261414 -902
rect 261954 680614 262574 711002
rect 271954 710598 272574 711590
rect 271954 710362 271986 710598
rect 272222 710362 272306 710598
rect 272542 710362 272574 710598
rect 271954 710278 272574 710362
rect 271954 710042 271986 710278
rect 272222 710042 272306 710278
rect 272542 710042 272574 710278
rect 268234 708678 268854 709670
rect 268234 708442 268266 708678
rect 268502 708442 268586 708678
rect 268822 708442 268854 708678
rect 268234 708358 268854 708442
rect 268234 708122 268266 708358
rect 268502 708122 268586 708358
rect 268822 708122 268854 708358
rect 261954 680378 261986 680614
rect 262222 680378 262306 680614
rect 262542 680378 262574 680614
rect 261954 680294 262574 680378
rect 261954 680058 261986 680294
rect 262222 680058 262306 680294
rect 262542 680058 262574 680294
rect 261954 644614 262574 680058
rect 261954 644378 261986 644614
rect 262222 644378 262306 644614
rect 262542 644378 262574 644614
rect 261954 644294 262574 644378
rect 261954 644058 261986 644294
rect 262222 644058 262306 644294
rect 262542 644058 262574 644294
rect 261954 608614 262574 644058
rect 261954 608378 261986 608614
rect 262222 608378 262306 608614
rect 262542 608378 262574 608614
rect 261954 608294 262574 608378
rect 261954 608058 261986 608294
rect 262222 608058 262306 608294
rect 262542 608058 262574 608294
rect 261954 572614 262574 608058
rect 261954 572378 261986 572614
rect 262222 572378 262306 572614
rect 262542 572378 262574 572614
rect 261954 572294 262574 572378
rect 261954 572058 261986 572294
rect 262222 572058 262306 572294
rect 262542 572058 262574 572294
rect 261954 536614 262574 572058
rect 261954 536378 261986 536614
rect 262222 536378 262306 536614
rect 262542 536378 262574 536614
rect 261954 536294 262574 536378
rect 261954 536058 261986 536294
rect 262222 536058 262306 536294
rect 262542 536058 262574 536294
rect 261954 500614 262574 536058
rect 261954 500378 261986 500614
rect 262222 500378 262306 500614
rect 262542 500378 262574 500614
rect 261954 500294 262574 500378
rect 261954 500058 261986 500294
rect 262222 500058 262306 500294
rect 262542 500058 262574 500294
rect 261954 464614 262574 500058
rect 261954 464378 261986 464614
rect 262222 464378 262306 464614
rect 262542 464378 262574 464614
rect 261954 464294 262574 464378
rect 261954 464058 261986 464294
rect 262222 464058 262306 464294
rect 262542 464058 262574 464294
rect 261954 428614 262574 464058
rect 261954 428378 261986 428614
rect 262222 428378 262306 428614
rect 262542 428378 262574 428614
rect 261954 428294 262574 428378
rect 261954 428058 261986 428294
rect 262222 428058 262306 428294
rect 262542 428058 262574 428294
rect 261954 392614 262574 428058
rect 261954 392378 261986 392614
rect 262222 392378 262306 392614
rect 262542 392378 262574 392614
rect 261954 392294 262574 392378
rect 261954 392058 261986 392294
rect 262222 392058 262306 392294
rect 262542 392058 262574 392294
rect 261954 356614 262574 392058
rect 261954 356378 261986 356614
rect 262222 356378 262306 356614
rect 262542 356378 262574 356614
rect 261954 356294 262574 356378
rect 261954 356058 261986 356294
rect 262222 356058 262306 356294
rect 262542 356058 262574 356294
rect 261954 320614 262574 356058
rect 261954 320378 261986 320614
rect 262222 320378 262306 320614
rect 262542 320378 262574 320614
rect 261954 320294 262574 320378
rect 261954 320058 261986 320294
rect 262222 320058 262306 320294
rect 262542 320058 262574 320294
rect 261954 284614 262574 320058
rect 261954 284378 261986 284614
rect 262222 284378 262306 284614
rect 262542 284378 262574 284614
rect 261954 284294 262574 284378
rect 261954 284058 261986 284294
rect 262222 284058 262306 284294
rect 262542 284058 262574 284294
rect 261954 248614 262574 284058
rect 261954 248378 261986 248614
rect 262222 248378 262306 248614
rect 262542 248378 262574 248614
rect 261954 248294 262574 248378
rect 261954 248058 261986 248294
rect 262222 248058 262306 248294
rect 262542 248058 262574 248294
rect 261954 212614 262574 248058
rect 261954 212378 261986 212614
rect 262222 212378 262306 212614
rect 262542 212378 262574 212614
rect 261954 212294 262574 212378
rect 261954 212058 261986 212294
rect 262222 212058 262306 212294
rect 262542 212058 262574 212294
rect 261954 176614 262574 212058
rect 261954 176378 261986 176614
rect 262222 176378 262306 176614
rect 262542 176378 262574 176614
rect 261954 176294 262574 176378
rect 261954 176058 261986 176294
rect 262222 176058 262306 176294
rect 262542 176058 262574 176294
rect 261954 140614 262574 176058
rect 261954 140378 261986 140614
rect 262222 140378 262306 140614
rect 262542 140378 262574 140614
rect 261954 140294 262574 140378
rect 261954 140058 261986 140294
rect 262222 140058 262306 140294
rect 262542 140058 262574 140294
rect 261954 104614 262574 140058
rect 261954 104378 261986 104614
rect 262222 104378 262306 104614
rect 262542 104378 262574 104614
rect 261954 104294 262574 104378
rect 261954 104058 261986 104294
rect 262222 104058 262306 104294
rect 262542 104058 262574 104294
rect 261954 68614 262574 104058
rect 261954 68378 261986 68614
rect 262222 68378 262306 68614
rect 262542 68378 262574 68614
rect 261954 68294 262574 68378
rect 261954 68058 261986 68294
rect 262222 68058 262306 68294
rect 262542 68058 262574 68294
rect 261954 32614 262574 68058
rect 261954 32378 261986 32614
rect 262222 32378 262306 32614
rect 262542 32378 262574 32614
rect 261954 32294 262574 32378
rect 261954 32058 261986 32294
rect 262222 32058 262306 32294
rect 262542 32058 262574 32294
rect 258234 -5382 258266 -5146
rect 258502 -5382 258586 -5146
rect 258822 -5382 258854 -5146
rect 258234 -5466 258854 -5382
rect 258234 -5702 258266 -5466
rect 258502 -5702 258586 -5466
rect 258822 -5702 258854 -5466
rect 258234 -5734 258854 -5702
rect 251954 -6342 251986 -6106
rect 252222 -6342 252306 -6106
rect 252542 -6342 252574 -6106
rect 251954 -6426 252574 -6342
rect 251954 -6662 251986 -6426
rect 252222 -6662 252306 -6426
rect 252542 -6662 252574 -6426
rect 251954 -7654 252574 -6662
rect 261954 -7066 262574 32058
rect 264514 706758 265134 707750
rect 264514 706522 264546 706758
rect 264782 706522 264866 706758
rect 265102 706522 265134 706758
rect 264514 706438 265134 706522
rect 264514 706202 264546 706438
rect 264782 706202 264866 706438
rect 265102 706202 265134 706438
rect 264514 691174 265134 706202
rect 264514 690938 264546 691174
rect 264782 690938 264866 691174
rect 265102 690938 265134 691174
rect 264514 690854 265134 690938
rect 264514 690618 264546 690854
rect 264782 690618 264866 690854
rect 265102 690618 265134 690854
rect 264514 655174 265134 690618
rect 264514 654938 264546 655174
rect 264782 654938 264866 655174
rect 265102 654938 265134 655174
rect 264514 654854 265134 654938
rect 264514 654618 264546 654854
rect 264782 654618 264866 654854
rect 265102 654618 265134 654854
rect 264514 619174 265134 654618
rect 264514 618938 264546 619174
rect 264782 618938 264866 619174
rect 265102 618938 265134 619174
rect 264514 618854 265134 618938
rect 264514 618618 264546 618854
rect 264782 618618 264866 618854
rect 265102 618618 265134 618854
rect 264514 583174 265134 618618
rect 264514 582938 264546 583174
rect 264782 582938 264866 583174
rect 265102 582938 265134 583174
rect 264514 582854 265134 582938
rect 264514 582618 264546 582854
rect 264782 582618 264866 582854
rect 265102 582618 265134 582854
rect 264514 547174 265134 582618
rect 264514 546938 264546 547174
rect 264782 546938 264866 547174
rect 265102 546938 265134 547174
rect 264514 546854 265134 546938
rect 264514 546618 264546 546854
rect 264782 546618 264866 546854
rect 265102 546618 265134 546854
rect 264514 511174 265134 546618
rect 264514 510938 264546 511174
rect 264782 510938 264866 511174
rect 265102 510938 265134 511174
rect 264514 510854 265134 510938
rect 264514 510618 264546 510854
rect 264782 510618 264866 510854
rect 265102 510618 265134 510854
rect 264514 475174 265134 510618
rect 264514 474938 264546 475174
rect 264782 474938 264866 475174
rect 265102 474938 265134 475174
rect 264514 474854 265134 474938
rect 264514 474618 264546 474854
rect 264782 474618 264866 474854
rect 265102 474618 265134 474854
rect 264514 439174 265134 474618
rect 264514 438938 264546 439174
rect 264782 438938 264866 439174
rect 265102 438938 265134 439174
rect 264514 438854 265134 438938
rect 264514 438618 264546 438854
rect 264782 438618 264866 438854
rect 265102 438618 265134 438854
rect 264514 403174 265134 438618
rect 264514 402938 264546 403174
rect 264782 402938 264866 403174
rect 265102 402938 265134 403174
rect 264514 402854 265134 402938
rect 264514 402618 264546 402854
rect 264782 402618 264866 402854
rect 265102 402618 265134 402854
rect 264514 367174 265134 402618
rect 264514 366938 264546 367174
rect 264782 366938 264866 367174
rect 265102 366938 265134 367174
rect 264514 366854 265134 366938
rect 264514 366618 264546 366854
rect 264782 366618 264866 366854
rect 265102 366618 265134 366854
rect 264514 331174 265134 366618
rect 264514 330938 264546 331174
rect 264782 330938 264866 331174
rect 265102 330938 265134 331174
rect 264514 330854 265134 330938
rect 264514 330618 264546 330854
rect 264782 330618 264866 330854
rect 265102 330618 265134 330854
rect 264514 295174 265134 330618
rect 264514 294938 264546 295174
rect 264782 294938 264866 295174
rect 265102 294938 265134 295174
rect 264514 294854 265134 294938
rect 264514 294618 264546 294854
rect 264782 294618 264866 294854
rect 265102 294618 265134 294854
rect 264514 259174 265134 294618
rect 264514 258938 264546 259174
rect 264782 258938 264866 259174
rect 265102 258938 265134 259174
rect 264514 258854 265134 258938
rect 264514 258618 264546 258854
rect 264782 258618 264866 258854
rect 265102 258618 265134 258854
rect 264514 223174 265134 258618
rect 264514 222938 264546 223174
rect 264782 222938 264866 223174
rect 265102 222938 265134 223174
rect 264514 222854 265134 222938
rect 264514 222618 264546 222854
rect 264782 222618 264866 222854
rect 265102 222618 265134 222854
rect 264514 187174 265134 222618
rect 264514 186938 264546 187174
rect 264782 186938 264866 187174
rect 265102 186938 265134 187174
rect 264514 186854 265134 186938
rect 264514 186618 264546 186854
rect 264782 186618 264866 186854
rect 265102 186618 265134 186854
rect 264514 151174 265134 186618
rect 264514 150938 264546 151174
rect 264782 150938 264866 151174
rect 265102 150938 265134 151174
rect 264514 150854 265134 150938
rect 264514 150618 264546 150854
rect 264782 150618 264866 150854
rect 265102 150618 265134 150854
rect 264514 115174 265134 150618
rect 264514 114938 264546 115174
rect 264782 114938 264866 115174
rect 265102 114938 265134 115174
rect 264514 114854 265134 114938
rect 264514 114618 264546 114854
rect 264782 114618 264866 114854
rect 265102 114618 265134 114854
rect 264514 79174 265134 114618
rect 264514 78938 264546 79174
rect 264782 78938 264866 79174
rect 265102 78938 265134 79174
rect 264514 78854 265134 78938
rect 264514 78618 264546 78854
rect 264782 78618 264866 78854
rect 265102 78618 265134 78854
rect 264514 43174 265134 78618
rect 264514 42938 264546 43174
rect 264782 42938 264866 43174
rect 265102 42938 265134 43174
rect 264514 42854 265134 42938
rect 264514 42618 264546 42854
rect 264782 42618 264866 42854
rect 265102 42618 265134 42854
rect 264514 7174 265134 42618
rect 264514 6938 264546 7174
rect 264782 6938 264866 7174
rect 265102 6938 265134 7174
rect 264514 6854 265134 6938
rect 264514 6618 264546 6854
rect 264782 6618 264866 6854
rect 265102 6618 265134 6854
rect 264514 -2266 265134 6618
rect 264514 -2502 264546 -2266
rect 264782 -2502 264866 -2266
rect 265102 -2502 265134 -2266
rect 264514 -2586 265134 -2502
rect 264514 -2822 264546 -2586
rect 264782 -2822 264866 -2586
rect 265102 -2822 265134 -2586
rect 264514 -3814 265134 -2822
rect 268234 694894 268854 708122
rect 268234 694658 268266 694894
rect 268502 694658 268586 694894
rect 268822 694658 268854 694894
rect 268234 694574 268854 694658
rect 268234 694338 268266 694574
rect 268502 694338 268586 694574
rect 268822 694338 268854 694574
rect 268234 658894 268854 694338
rect 268234 658658 268266 658894
rect 268502 658658 268586 658894
rect 268822 658658 268854 658894
rect 268234 658574 268854 658658
rect 268234 658338 268266 658574
rect 268502 658338 268586 658574
rect 268822 658338 268854 658574
rect 268234 622894 268854 658338
rect 268234 622658 268266 622894
rect 268502 622658 268586 622894
rect 268822 622658 268854 622894
rect 268234 622574 268854 622658
rect 268234 622338 268266 622574
rect 268502 622338 268586 622574
rect 268822 622338 268854 622574
rect 268234 586894 268854 622338
rect 268234 586658 268266 586894
rect 268502 586658 268586 586894
rect 268822 586658 268854 586894
rect 268234 586574 268854 586658
rect 268234 586338 268266 586574
rect 268502 586338 268586 586574
rect 268822 586338 268854 586574
rect 268234 550894 268854 586338
rect 268234 550658 268266 550894
rect 268502 550658 268586 550894
rect 268822 550658 268854 550894
rect 268234 550574 268854 550658
rect 268234 550338 268266 550574
rect 268502 550338 268586 550574
rect 268822 550338 268854 550574
rect 268234 514894 268854 550338
rect 268234 514658 268266 514894
rect 268502 514658 268586 514894
rect 268822 514658 268854 514894
rect 268234 514574 268854 514658
rect 268234 514338 268266 514574
rect 268502 514338 268586 514574
rect 268822 514338 268854 514574
rect 268234 478894 268854 514338
rect 268234 478658 268266 478894
rect 268502 478658 268586 478894
rect 268822 478658 268854 478894
rect 268234 478574 268854 478658
rect 268234 478338 268266 478574
rect 268502 478338 268586 478574
rect 268822 478338 268854 478574
rect 268234 442894 268854 478338
rect 268234 442658 268266 442894
rect 268502 442658 268586 442894
rect 268822 442658 268854 442894
rect 268234 442574 268854 442658
rect 268234 442338 268266 442574
rect 268502 442338 268586 442574
rect 268822 442338 268854 442574
rect 268234 406894 268854 442338
rect 268234 406658 268266 406894
rect 268502 406658 268586 406894
rect 268822 406658 268854 406894
rect 268234 406574 268854 406658
rect 268234 406338 268266 406574
rect 268502 406338 268586 406574
rect 268822 406338 268854 406574
rect 268234 370894 268854 406338
rect 268234 370658 268266 370894
rect 268502 370658 268586 370894
rect 268822 370658 268854 370894
rect 268234 370574 268854 370658
rect 268234 370338 268266 370574
rect 268502 370338 268586 370574
rect 268822 370338 268854 370574
rect 268234 334894 268854 370338
rect 268234 334658 268266 334894
rect 268502 334658 268586 334894
rect 268822 334658 268854 334894
rect 268234 334574 268854 334658
rect 268234 334338 268266 334574
rect 268502 334338 268586 334574
rect 268822 334338 268854 334574
rect 268234 298894 268854 334338
rect 268234 298658 268266 298894
rect 268502 298658 268586 298894
rect 268822 298658 268854 298894
rect 268234 298574 268854 298658
rect 268234 298338 268266 298574
rect 268502 298338 268586 298574
rect 268822 298338 268854 298574
rect 268234 262894 268854 298338
rect 268234 262658 268266 262894
rect 268502 262658 268586 262894
rect 268822 262658 268854 262894
rect 268234 262574 268854 262658
rect 268234 262338 268266 262574
rect 268502 262338 268586 262574
rect 268822 262338 268854 262574
rect 268234 226894 268854 262338
rect 268234 226658 268266 226894
rect 268502 226658 268586 226894
rect 268822 226658 268854 226894
rect 268234 226574 268854 226658
rect 268234 226338 268266 226574
rect 268502 226338 268586 226574
rect 268822 226338 268854 226574
rect 268234 190894 268854 226338
rect 268234 190658 268266 190894
rect 268502 190658 268586 190894
rect 268822 190658 268854 190894
rect 268234 190574 268854 190658
rect 268234 190338 268266 190574
rect 268502 190338 268586 190574
rect 268822 190338 268854 190574
rect 268234 154894 268854 190338
rect 268234 154658 268266 154894
rect 268502 154658 268586 154894
rect 268822 154658 268854 154894
rect 268234 154574 268854 154658
rect 268234 154338 268266 154574
rect 268502 154338 268586 154574
rect 268822 154338 268854 154574
rect 268234 118894 268854 154338
rect 268234 118658 268266 118894
rect 268502 118658 268586 118894
rect 268822 118658 268854 118894
rect 268234 118574 268854 118658
rect 268234 118338 268266 118574
rect 268502 118338 268586 118574
rect 268822 118338 268854 118574
rect 268234 82894 268854 118338
rect 268234 82658 268266 82894
rect 268502 82658 268586 82894
rect 268822 82658 268854 82894
rect 268234 82574 268854 82658
rect 268234 82338 268266 82574
rect 268502 82338 268586 82574
rect 268822 82338 268854 82574
rect 268234 46894 268854 82338
rect 268234 46658 268266 46894
rect 268502 46658 268586 46894
rect 268822 46658 268854 46894
rect 268234 46574 268854 46658
rect 268234 46338 268266 46574
rect 268502 46338 268586 46574
rect 268822 46338 268854 46574
rect 268234 10894 268854 46338
rect 268234 10658 268266 10894
rect 268502 10658 268586 10894
rect 268822 10658 268854 10894
rect 268234 10574 268854 10658
rect 268234 10338 268266 10574
rect 268502 10338 268586 10574
rect 268822 10338 268854 10574
rect 268234 -4186 268854 10338
rect 270794 705798 271414 705830
rect 270794 705562 270826 705798
rect 271062 705562 271146 705798
rect 271382 705562 271414 705798
rect 270794 705478 271414 705562
rect 270794 705242 270826 705478
rect 271062 705242 271146 705478
rect 271382 705242 271414 705478
rect 270794 669454 271414 705242
rect 270794 669218 270826 669454
rect 271062 669218 271146 669454
rect 271382 669218 271414 669454
rect 270794 669134 271414 669218
rect 270794 668898 270826 669134
rect 271062 668898 271146 669134
rect 271382 668898 271414 669134
rect 270794 633454 271414 668898
rect 270794 633218 270826 633454
rect 271062 633218 271146 633454
rect 271382 633218 271414 633454
rect 270794 633134 271414 633218
rect 270794 632898 270826 633134
rect 271062 632898 271146 633134
rect 271382 632898 271414 633134
rect 270794 597454 271414 632898
rect 270794 597218 270826 597454
rect 271062 597218 271146 597454
rect 271382 597218 271414 597454
rect 270794 597134 271414 597218
rect 270794 596898 270826 597134
rect 271062 596898 271146 597134
rect 271382 596898 271414 597134
rect 270794 561454 271414 596898
rect 270794 561218 270826 561454
rect 271062 561218 271146 561454
rect 271382 561218 271414 561454
rect 270794 561134 271414 561218
rect 270794 560898 270826 561134
rect 271062 560898 271146 561134
rect 271382 560898 271414 561134
rect 270794 525454 271414 560898
rect 270794 525218 270826 525454
rect 271062 525218 271146 525454
rect 271382 525218 271414 525454
rect 270794 525134 271414 525218
rect 270794 524898 270826 525134
rect 271062 524898 271146 525134
rect 271382 524898 271414 525134
rect 270794 489454 271414 524898
rect 270794 489218 270826 489454
rect 271062 489218 271146 489454
rect 271382 489218 271414 489454
rect 270794 489134 271414 489218
rect 270794 488898 270826 489134
rect 271062 488898 271146 489134
rect 271382 488898 271414 489134
rect 270794 453454 271414 488898
rect 270794 453218 270826 453454
rect 271062 453218 271146 453454
rect 271382 453218 271414 453454
rect 270794 453134 271414 453218
rect 270794 452898 270826 453134
rect 271062 452898 271146 453134
rect 271382 452898 271414 453134
rect 270794 417454 271414 452898
rect 270794 417218 270826 417454
rect 271062 417218 271146 417454
rect 271382 417218 271414 417454
rect 270794 417134 271414 417218
rect 270794 416898 270826 417134
rect 271062 416898 271146 417134
rect 271382 416898 271414 417134
rect 270794 381454 271414 416898
rect 270794 381218 270826 381454
rect 271062 381218 271146 381454
rect 271382 381218 271414 381454
rect 270794 381134 271414 381218
rect 270794 380898 270826 381134
rect 271062 380898 271146 381134
rect 271382 380898 271414 381134
rect 270794 345454 271414 380898
rect 270794 345218 270826 345454
rect 271062 345218 271146 345454
rect 271382 345218 271414 345454
rect 270794 345134 271414 345218
rect 270794 344898 270826 345134
rect 271062 344898 271146 345134
rect 271382 344898 271414 345134
rect 270794 309454 271414 344898
rect 270794 309218 270826 309454
rect 271062 309218 271146 309454
rect 271382 309218 271414 309454
rect 270794 309134 271414 309218
rect 270794 308898 270826 309134
rect 271062 308898 271146 309134
rect 271382 308898 271414 309134
rect 270794 273454 271414 308898
rect 270794 273218 270826 273454
rect 271062 273218 271146 273454
rect 271382 273218 271414 273454
rect 270794 273134 271414 273218
rect 270794 272898 270826 273134
rect 271062 272898 271146 273134
rect 271382 272898 271414 273134
rect 270794 237454 271414 272898
rect 270794 237218 270826 237454
rect 271062 237218 271146 237454
rect 271382 237218 271414 237454
rect 270794 237134 271414 237218
rect 270794 236898 270826 237134
rect 271062 236898 271146 237134
rect 271382 236898 271414 237134
rect 270794 201454 271414 236898
rect 270794 201218 270826 201454
rect 271062 201218 271146 201454
rect 271382 201218 271414 201454
rect 270794 201134 271414 201218
rect 270794 200898 270826 201134
rect 271062 200898 271146 201134
rect 271382 200898 271414 201134
rect 270794 165454 271414 200898
rect 270794 165218 270826 165454
rect 271062 165218 271146 165454
rect 271382 165218 271414 165454
rect 270794 165134 271414 165218
rect 270794 164898 270826 165134
rect 271062 164898 271146 165134
rect 271382 164898 271414 165134
rect 270794 129454 271414 164898
rect 270794 129218 270826 129454
rect 271062 129218 271146 129454
rect 271382 129218 271414 129454
rect 270794 129134 271414 129218
rect 270794 128898 270826 129134
rect 271062 128898 271146 129134
rect 271382 128898 271414 129134
rect 270794 93454 271414 128898
rect 270794 93218 270826 93454
rect 271062 93218 271146 93454
rect 271382 93218 271414 93454
rect 270794 93134 271414 93218
rect 270794 92898 270826 93134
rect 271062 92898 271146 93134
rect 271382 92898 271414 93134
rect 270794 57454 271414 92898
rect 270794 57218 270826 57454
rect 271062 57218 271146 57454
rect 271382 57218 271414 57454
rect 270794 57134 271414 57218
rect 270794 56898 270826 57134
rect 271062 56898 271146 57134
rect 271382 56898 271414 57134
rect 270794 21454 271414 56898
rect 270794 21218 270826 21454
rect 271062 21218 271146 21454
rect 271382 21218 271414 21454
rect 270794 21134 271414 21218
rect 270794 20898 270826 21134
rect 271062 20898 271146 21134
rect 271382 20898 271414 21134
rect 270794 -1306 271414 20898
rect 270794 -1542 270826 -1306
rect 271062 -1542 271146 -1306
rect 271382 -1542 271414 -1306
rect 270794 -1626 271414 -1542
rect 270794 -1862 270826 -1626
rect 271062 -1862 271146 -1626
rect 271382 -1862 271414 -1626
rect 270794 -1894 271414 -1862
rect 271954 698614 272574 710042
rect 281954 711558 282574 711590
rect 281954 711322 281986 711558
rect 282222 711322 282306 711558
rect 282542 711322 282574 711558
rect 281954 711238 282574 711322
rect 281954 711002 281986 711238
rect 282222 711002 282306 711238
rect 282542 711002 282574 711238
rect 278234 709638 278854 709670
rect 278234 709402 278266 709638
rect 278502 709402 278586 709638
rect 278822 709402 278854 709638
rect 278234 709318 278854 709402
rect 278234 709082 278266 709318
rect 278502 709082 278586 709318
rect 278822 709082 278854 709318
rect 271954 698378 271986 698614
rect 272222 698378 272306 698614
rect 272542 698378 272574 698614
rect 271954 698294 272574 698378
rect 271954 698058 271986 698294
rect 272222 698058 272306 698294
rect 272542 698058 272574 698294
rect 271954 662614 272574 698058
rect 271954 662378 271986 662614
rect 272222 662378 272306 662614
rect 272542 662378 272574 662614
rect 271954 662294 272574 662378
rect 271954 662058 271986 662294
rect 272222 662058 272306 662294
rect 272542 662058 272574 662294
rect 271954 626614 272574 662058
rect 271954 626378 271986 626614
rect 272222 626378 272306 626614
rect 272542 626378 272574 626614
rect 271954 626294 272574 626378
rect 271954 626058 271986 626294
rect 272222 626058 272306 626294
rect 272542 626058 272574 626294
rect 271954 590614 272574 626058
rect 271954 590378 271986 590614
rect 272222 590378 272306 590614
rect 272542 590378 272574 590614
rect 271954 590294 272574 590378
rect 271954 590058 271986 590294
rect 272222 590058 272306 590294
rect 272542 590058 272574 590294
rect 271954 554614 272574 590058
rect 271954 554378 271986 554614
rect 272222 554378 272306 554614
rect 272542 554378 272574 554614
rect 271954 554294 272574 554378
rect 271954 554058 271986 554294
rect 272222 554058 272306 554294
rect 272542 554058 272574 554294
rect 271954 518614 272574 554058
rect 271954 518378 271986 518614
rect 272222 518378 272306 518614
rect 272542 518378 272574 518614
rect 271954 518294 272574 518378
rect 271954 518058 271986 518294
rect 272222 518058 272306 518294
rect 272542 518058 272574 518294
rect 271954 482614 272574 518058
rect 271954 482378 271986 482614
rect 272222 482378 272306 482614
rect 272542 482378 272574 482614
rect 271954 482294 272574 482378
rect 271954 482058 271986 482294
rect 272222 482058 272306 482294
rect 272542 482058 272574 482294
rect 271954 446614 272574 482058
rect 271954 446378 271986 446614
rect 272222 446378 272306 446614
rect 272542 446378 272574 446614
rect 271954 446294 272574 446378
rect 271954 446058 271986 446294
rect 272222 446058 272306 446294
rect 272542 446058 272574 446294
rect 271954 410614 272574 446058
rect 271954 410378 271986 410614
rect 272222 410378 272306 410614
rect 272542 410378 272574 410614
rect 271954 410294 272574 410378
rect 271954 410058 271986 410294
rect 272222 410058 272306 410294
rect 272542 410058 272574 410294
rect 271954 374614 272574 410058
rect 271954 374378 271986 374614
rect 272222 374378 272306 374614
rect 272542 374378 272574 374614
rect 271954 374294 272574 374378
rect 271954 374058 271986 374294
rect 272222 374058 272306 374294
rect 272542 374058 272574 374294
rect 271954 338614 272574 374058
rect 271954 338378 271986 338614
rect 272222 338378 272306 338614
rect 272542 338378 272574 338614
rect 271954 338294 272574 338378
rect 271954 338058 271986 338294
rect 272222 338058 272306 338294
rect 272542 338058 272574 338294
rect 271954 302614 272574 338058
rect 271954 302378 271986 302614
rect 272222 302378 272306 302614
rect 272542 302378 272574 302614
rect 271954 302294 272574 302378
rect 271954 302058 271986 302294
rect 272222 302058 272306 302294
rect 272542 302058 272574 302294
rect 271954 266614 272574 302058
rect 271954 266378 271986 266614
rect 272222 266378 272306 266614
rect 272542 266378 272574 266614
rect 271954 266294 272574 266378
rect 271954 266058 271986 266294
rect 272222 266058 272306 266294
rect 272542 266058 272574 266294
rect 271954 230614 272574 266058
rect 271954 230378 271986 230614
rect 272222 230378 272306 230614
rect 272542 230378 272574 230614
rect 271954 230294 272574 230378
rect 271954 230058 271986 230294
rect 272222 230058 272306 230294
rect 272542 230058 272574 230294
rect 271954 194614 272574 230058
rect 271954 194378 271986 194614
rect 272222 194378 272306 194614
rect 272542 194378 272574 194614
rect 271954 194294 272574 194378
rect 271954 194058 271986 194294
rect 272222 194058 272306 194294
rect 272542 194058 272574 194294
rect 271954 158614 272574 194058
rect 271954 158378 271986 158614
rect 272222 158378 272306 158614
rect 272542 158378 272574 158614
rect 271954 158294 272574 158378
rect 271954 158058 271986 158294
rect 272222 158058 272306 158294
rect 272542 158058 272574 158294
rect 271954 122614 272574 158058
rect 271954 122378 271986 122614
rect 272222 122378 272306 122614
rect 272542 122378 272574 122614
rect 271954 122294 272574 122378
rect 271954 122058 271986 122294
rect 272222 122058 272306 122294
rect 272542 122058 272574 122294
rect 271954 86614 272574 122058
rect 271954 86378 271986 86614
rect 272222 86378 272306 86614
rect 272542 86378 272574 86614
rect 271954 86294 272574 86378
rect 271954 86058 271986 86294
rect 272222 86058 272306 86294
rect 272542 86058 272574 86294
rect 271954 50614 272574 86058
rect 271954 50378 271986 50614
rect 272222 50378 272306 50614
rect 272542 50378 272574 50614
rect 271954 50294 272574 50378
rect 271954 50058 271986 50294
rect 272222 50058 272306 50294
rect 272542 50058 272574 50294
rect 271954 14614 272574 50058
rect 271954 14378 271986 14614
rect 272222 14378 272306 14614
rect 272542 14378 272574 14614
rect 271954 14294 272574 14378
rect 271954 14058 271986 14294
rect 272222 14058 272306 14294
rect 272542 14058 272574 14294
rect 268234 -4422 268266 -4186
rect 268502 -4422 268586 -4186
rect 268822 -4422 268854 -4186
rect 268234 -4506 268854 -4422
rect 268234 -4742 268266 -4506
rect 268502 -4742 268586 -4506
rect 268822 -4742 268854 -4506
rect 268234 -5734 268854 -4742
rect 261954 -7302 261986 -7066
rect 262222 -7302 262306 -7066
rect 262542 -7302 262574 -7066
rect 261954 -7386 262574 -7302
rect 261954 -7622 261986 -7386
rect 262222 -7622 262306 -7386
rect 262542 -7622 262574 -7386
rect 261954 -7654 262574 -7622
rect 271954 -6106 272574 14058
rect 274514 707718 275134 707750
rect 274514 707482 274546 707718
rect 274782 707482 274866 707718
rect 275102 707482 275134 707718
rect 274514 707398 275134 707482
rect 274514 707162 274546 707398
rect 274782 707162 274866 707398
rect 275102 707162 275134 707398
rect 274514 673174 275134 707162
rect 274514 672938 274546 673174
rect 274782 672938 274866 673174
rect 275102 672938 275134 673174
rect 274514 672854 275134 672938
rect 274514 672618 274546 672854
rect 274782 672618 274866 672854
rect 275102 672618 275134 672854
rect 274514 637174 275134 672618
rect 274514 636938 274546 637174
rect 274782 636938 274866 637174
rect 275102 636938 275134 637174
rect 274514 636854 275134 636938
rect 274514 636618 274546 636854
rect 274782 636618 274866 636854
rect 275102 636618 275134 636854
rect 274514 601174 275134 636618
rect 274514 600938 274546 601174
rect 274782 600938 274866 601174
rect 275102 600938 275134 601174
rect 274514 600854 275134 600938
rect 274514 600618 274546 600854
rect 274782 600618 274866 600854
rect 275102 600618 275134 600854
rect 274514 565174 275134 600618
rect 274514 564938 274546 565174
rect 274782 564938 274866 565174
rect 275102 564938 275134 565174
rect 274514 564854 275134 564938
rect 274514 564618 274546 564854
rect 274782 564618 274866 564854
rect 275102 564618 275134 564854
rect 274514 529174 275134 564618
rect 274514 528938 274546 529174
rect 274782 528938 274866 529174
rect 275102 528938 275134 529174
rect 274514 528854 275134 528938
rect 274514 528618 274546 528854
rect 274782 528618 274866 528854
rect 275102 528618 275134 528854
rect 274514 493174 275134 528618
rect 274514 492938 274546 493174
rect 274782 492938 274866 493174
rect 275102 492938 275134 493174
rect 274514 492854 275134 492938
rect 274514 492618 274546 492854
rect 274782 492618 274866 492854
rect 275102 492618 275134 492854
rect 274514 457174 275134 492618
rect 274514 456938 274546 457174
rect 274782 456938 274866 457174
rect 275102 456938 275134 457174
rect 274514 456854 275134 456938
rect 274514 456618 274546 456854
rect 274782 456618 274866 456854
rect 275102 456618 275134 456854
rect 274514 421174 275134 456618
rect 274514 420938 274546 421174
rect 274782 420938 274866 421174
rect 275102 420938 275134 421174
rect 274514 420854 275134 420938
rect 274514 420618 274546 420854
rect 274782 420618 274866 420854
rect 275102 420618 275134 420854
rect 274514 385174 275134 420618
rect 274514 384938 274546 385174
rect 274782 384938 274866 385174
rect 275102 384938 275134 385174
rect 274514 384854 275134 384938
rect 274514 384618 274546 384854
rect 274782 384618 274866 384854
rect 275102 384618 275134 384854
rect 274514 349174 275134 384618
rect 274514 348938 274546 349174
rect 274782 348938 274866 349174
rect 275102 348938 275134 349174
rect 274514 348854 275134 348938
rect 274514 348618 274546 348854
rect 274782 348618 274866 348854
rect 275102 348618 275134 348854
rect 274514 313174 275134 348618
rect 274514 312938 274546 313174
rect 274782 312938 274866 313174
rect 275102 312938 275134 313174
rect 274514 312854 275134 312938
rect 274514 312618 274546 312854
rect 274782 312618 274866 312854
rect 275102 312618 275134 312854
rect 274514 277174 275134 312618
rect 274514 276938 274546 277174
rect 274782 276938 274866 277174
rect 275102 276938 275134 277174
rect 274514 276854 275134 276938
rect 274514 276618 274546 276854
rect 274782 276618 274866 276854
rect 275102 276618 275134 276854
rect 274514 241174 275134 276618
rect 274514 240938 274546 241174
rect 274782 240938 274866 241174
rect 275102 240938 275134 241174
rect 274514 240854 275134 240938
rect 274514 240618 274546 240854
rect 274782 240618 274866 240854
rect 275102 240618 275134 240854
rect 274514 205174 275134 240618
rect 274514 204938 274546 205174
rect 274782 204938 274866 205174
rect 275102 204938 275134 205174
rect 274514 204854 275134 204938
rect 274514 204618 274546 204854
rect 274782 204618 274866 204854
rect 275102 204618 275134 204854
rect 274514 169174 275134 204618
rect 274514 168938 274546 169174
rect 274782 168938 274866 169174
rect 275102 168938 275134 169174
rect 274514 168854 275134 168938
rect 274514 168618 274546 168854
rect 274782 168618 274866 168854
rect 275102 168618 275134 168854
rect 274514 133174 275134 168618
rect 274514 132938 274546 133174
rect 274782 132938 274866 133174
rect 275102 132938 275134 133174
rect 274514 132854 275134 132938
rect 274514 132618 274546 132854
rect 274782 132618 274866 132854
rect 275102 132618 275134 132854
rect 274514 97174 275134 132618
rect 274514 96938 274546 97174
rect 274782 96938 274866 97174
rect 275102 96938 275134 97174
rect 274514 96854 275134 96938
rect 274514 96618 274546 96854
rect 274782 96618 274866 96854
rect 275102 96618 275134 96854
rect 274514 61174 275134 96618
rect 274514 60938 274546 61174
rect 274782 60938 274866 61174
rect 275102 60938 275134 61174
rect 274514 60854 275134 60938
rect 274514 60618 274546 60854
rect 274782 60618 274866 60854
rect 275102 60618 275134 60854
rect 274514 25174 275134 60618
rect 274514 24938 274546 25174
rect 274782 24938 274866 25174
rect 275102 24938 275134 25174
rect 274514 24854 275134 24938
rect 274514 24618 274546 24854
rect 274782 24618 274866 24854
rect 275102 24618 275134 24854
rect 274514 -3226 275134 24618
rect 274514 -3462 274546 -3226
rect 274782 -3462 274866 -3226
rect 275102 -3462 275134 -3226
rect 274514 -3546 275134 -3462
rect 274514 -3782 274546 -3546
rect 274782 -3782 274866 -3546
rect 275102 -3782 275134 -3546
rect 274514 -3814 275134 -3782
rect 278234 676894 278854 709082
rect 278234 676658 278266 676894
rect 278502 676658 278586 676894
rect 278822 676658 278854 676894
rect 278234 676574 278854 676658
rect 278234 676338 278266 676574
rect 278502 676338 278586 676574
rect 278822 676338 278854 676574
rect 278234 640894 278854 676338
rect 278234 640658 278266 640894
rect 278502 640658 278586 640894
rect 278822 640658 278854 640894
rect 278234 640574 278854 640658
rect 278234 640338 278266 640574
rect 278502 640338 278586 640574
rect 278822 640338 278854 640574
rect 278234 604894 278854 640338
rect 278234 604658 278266 604894
rect 278502 604658 278586 604894
rect 278822 604658 278854 604894
rect 278234 604574 278854 604658
rect 278234 604338 278266 604574
rect 278502 604338 278586 604574
rect 278822 604338 278854 604574
rect 278234 568894 278854 604338
rect 278234 568658 278266 568894
rect 278502 568658 278586 568894
rect 278822 568658 278854 568894
rect 278234 568574 278854 568658
rect 278234 568338 278266 568574
rect 278502 568338 278586 568574
rect 278822 568338 278854 568574
rect 278234 532894 278854 568338
rect 278234 532658 278266 532894
rect 278502 532658 278586 532894
rect 278822 532658 278854 532894
rect 278234 532574 278854 532658
rect 278234 532338 278266 532574
rect 278502 532338 278586 532574
rect 278822 532338 278854 532574
rect 278234 496894 278854 532338
rect 278234 496658 278266 496894
rect 278502 496658 278586 496894
rect 278822 496658 278854 496894
rect 278234 496574 278854 496658
rect 278234 496338 278266 496574
rect 278502 496338 278586 496574
rect 278822 496338 278854 496574
rect 278234 460894 278854 496338
rect 278234 460658 278266 460894
rect 278502 460658 278586 460894
rect 278822 460658 278854 460894
rect 278234 460574 278854 460658
rect 278234 460338 278266 460574
rect 278502 460338 278586 460574
rect 278822 460338 278854 460574
rect 278234 424894 278854 460338
rect 278234 424658 278266 424894
rect 278502 424658 278586 424894
rect 278822 424658 278854 424894
rect 278234 424574 278854 424658
rect 278234 424338 278266 424574
rect 278502 424338 278586 424574
rect 278822 424338 278854 424574
rect 278234 388894 278854 424338
rect 278234 388658 278266 388894
rect 278502 388658 278586 388894
rect 278822 388658 278854 388894
rect 278234 388574 278854 388658
rect 278234 388338 278266 388574
rect 278502 388338 278586 388574
rect 278822 388338 278854 388574
rect 278234 352894 278854 388338
rect 278234 352658 278266 352894
rect 278502 352658 278586 352894
rect 278822 352658 278854 352894
rect 278234 352574 278854 352658
rect 278234 352338 278266 352574
rect 278502 352338 278586 352574
rect 278822 352338 278854 352574
rect 278234 316894 278854 352338
rect 278234 316658 278266 316894
rect 278502 316658 278586 316894
rect 278822 316658 278854 316894
rect 278234 316574 278854 316658
rect 278234 316338 278266 316574
rect 278502 316338 278586 316574
rect 278822 316338 278854 316574
rect 278234 280894 278854 316338
rect 278234 280658 278266 280894
rect 278502 280658 278586 280894
rect 278822 280658 278854 280894
rect 278234 280574 278854 280658
rect 278234 280338 278266 280574
rect 278502 280338 278586 280574
rect 278822 280338 278854 280574
rect 278234 244894 278854 280338
rect 278234 244658 278266 244894
rect 278502 244658 278586 244894
rect 278822 244658 278854 244894
rect 278234 244574 278854 244658
rect 278234 244338 278266 244574
rect 278502 244338 278586 244574
rect 278822 244338 278854 244574
rect 278234 208894 278854 244338
rect 278234 208658 278266 208894
rect 278502 208658 278586 208894
rect 278822 208658 278854 208894
rect 278234 208574 278854 208658
rect 278234 208338 278266 208574
rect 278502 208338 278586 208574
rect 278822 208338 278854 208574
rect 278234 172894 278854 208338
rect 278234 172658 278266 172894
rect 278502 172658 278586 172894
rect 278822 172658 278854 172894
rect 278234 172574 278854 172658
rect 278234 172338 278266 172574
rect 278502 172338 278586 172574
rect 278822 172338 278854 172574
rect 278234 136894 278854 172338
rect 278234 136658 278266 136894
rect 278502 136658 278586 136894
rect 278822 136658 278854 136894
rect 278234 136574 278854 136658
rect 278234 136338 278266 136574
rect 278502 136338 278586 136574
rect 278822 136338 278854 136574
rect 278234 100894 278854 136338
rect 278234 100658 278266 100894
rect 278502 100658 278586 100894
rect 278822 100658 278854 100894
rect 278234 100574 278854 100658
rect 278234 100338 278266 100574
rect 278502 100338 278586 100574
rect 278822 100338 278854 100574
rect 278234 64894 278854 100338
rect 278234 64658 278266 64894
rect 278502 64658 278586 64894
rect 278822 64658 278854 64894
rect 278234 64574 278854 64658
rect 278234 64338 278266 64574
rect 278502 64338 278586 64574
rect 278822 64338 278854 64574
rect 278234 28894 278854 64338
rect 278234 28658 278266 28894
rect 278502 28658 278586 28894
rect 278822 28658 278854 28894
rect 278234 28574 278854 28658
rect 278234 28338 278266 28574
rect 278502 28338 278586 28574
rect 278822 28338 278854 28574
rect 278234 -5146 278854 28338
rect 280794 704838 281414 705830
rect 280794 704602 280826 704838
rect 281062 704602 281146 704838
rect 281382 704602 281414 704838
rect 280794 704518 281414 704602
rect 280794 704282 280826 704518
rect 281062 704282 281146 704518
rect 281382 704282 281414 704518
rect 280794 687454 281414 704282
rect 280794 687218 280826 687454
rect 281062 687218 281146 687454
rect 281382 687218 281414 687454
rect 280794 687134 281414 687218
rect 280794 686898 280826 687134
rect 281062 686898 281146 687134
rect 281382 686898 281414 687134
rect 280794 651454 281414 686898
rect 280794 651218 280826 651454
rect 281062 651218 281146 651454
rect 281382 651218 281414 651454
rect 280794 651134 281414 651218
rect 280794 650898 280826 651134
rect 281062 650898 281146 651134
rect 281382 650898 281414 651134
rect 280794 615454 281414 650898
rect 280794 615218 280826 615454
rect 281062 615218 281146 615454
rect 281382 615218 281414 615454
rect 280794 615134 281414 615218
rect 280794 614898 280826 615134
rect 281062 614898 281146 615134
rect 281382 614898 281414 615134
rect 280794 579454 281414 614898
rect 280794 579218 280826 579454
rect 281062 579218 281146 579454
rect 281382 579218 281414 579454
rect 280794 579134 281414 579218
rect 280794 578898 280826 579134
rect 281062 578898 281146 579134
rect 281382 578898 281414 579134
rect 280794 543454 281414 578898
rect 280794 543218 280826 543454
rect 281062 543218 281146 543454
rect 281382 543218 281414 543454
rect 280794 543134 281414 543218
rect 280794 542898 280826 543134
rect 281062 542898 281146 543134
rect 281382 542898 281414 543134
rect 280794 507454 281414 542898
rect 280794 507218 280826 507454
rect 281062 507218 281146 507454
rect 281382 507218 281414 507454
rect 280794 507134 281414 507218
rect 280794 506898 280826 507134
rect 281062 506898 281146 507134
rect 281382 506898 281414 507134
rect 280794 471454 281414 506898
rect 280794 471218 280826 471454
rect 281062 471218 281146 471454
rect 281382 471218 281414 471454
rect 280794 471134 281414 471218
rect 280794 470898 280826 471134
rect 281062 470898 281146 471134
rect 281382 470898 281414 471134
rect 280794 435454 281414 470898
rect 280794 435218 280826 435454
rect 281062 435218 281146 435454
rect 281382 435218 281414 435454
rect 280794 435134 281414 435218
rect 280794 434898 280826 435134
rect 281062 434898 281146 435134
rect 281382 434898 281414 435134
rect 280794 399454 281414 434898
rect 280794 399218 280826 399454
rect 281062 399218 281146 399454
rect 281382 399218 281414 399454
rect 280794 399134 281414 399218
rect 280794 398898 280826 399134
rect 281062 398898 281146 399134
rect 281382 398898 281414 399134
rect 280794 363454 281414 398898
rect 280794 363218 280826 363454
rect 281062 363218 281146 363454
rect 281382 363218 281414 363454
rect 280794 363134 281414 363218
rect 280794 362898 280826 363134
rect 281062 362898 281146 363134
rect 281382 362898 281414 363134
rect 280794 327454 281414 362898
rect 280794 327218 280826 327454
rect 281062 327218 281146 327454
rect 281382 327218 281414 327454
rect 280794 327134 281414 327218
rect 280794 326898 280826 327134
rect 281062 326898 281146 327134
rect 281382 326898 281414 327134
rect 280794 291454 281414 326898
rect 280794 291218 280826 291454
rect 281062 291218 281146 291454
rect 281382 291218 281414 291454
rect 280794 291134 281414 291218
rect 280794 290898 280826 291134
rect 281062 290898 281146 291134
rect 281382 290898 281414 291134
rect 280794 255454 281414 290898
rect 280794 255218 280826 255454
rect 281062 255218 281146 255454
rect 281382 255218 281414 255454
rect 280794 255134 281414 255218
rect 280794 254898 280826 255134
rect 281062 254898 281146 255134
rect 281382 254898 281414 255134
rect 280794 219454 281414 254898
rect 280794 219218 280826 219454
rect 281062 219218 281146 219454
rect 281382 219218 281414 219454
rect 280794 219134 281414 219218
rect 280794 218898 280826 219134
rect 281062 218898 281146 219134
rect 281382 218898 281414 219134
rect 280794 183454 281414 218898
rect 280794 183218 280826 183454
rect 281062 183218 281146 183454
rect 281382 183218 281414 183454
rect 280794 183134 281414 183218
rect 280794 182898 280826 183134
rect 281062 182898 281146 183134
rect 281382 182898 281414 183134
rect 280794 147454 281414 182898
rect 280794 147218 280826 147454
rect 281062 147218 281146 147454
rect 281382 147218 281414 147454
rect 280794 147134 281414 147218
rect 280794 146898 280826 147134
rect 281062 146898 281146 147134
rect 281382 146898 281414 147134
rect 280794 111454 281414 146898
rect 280794 111218 280826 111454
rect 281062 111218 281146 111454
rect 281382 111218 281414 111454
rect 280794 111134 281414 111218
rect 280794 110898 280826 111134
rect 281062 110898 281146 111134
rect 281382 110898 281414 111134
rect 280794 75454 281414 110898
rect 280794 75218 280826 75454
rect 281062 75218 281146 75454
rect 281382 75218 281414 75454
rect 280794 75134 281414 75218
rect 280794 74898 280826 75134
rect 281062 74898 281146 75134
rect 281382 74898 281414 75134
rect 280794 39454 281414 74898
rect 280794 39218 280826 39454
rect 281062 39218 281146 39454
rect 281382 39218 281414 39454
rect 280794 39134 281414 39218
rect 280794 38898 280826 39134
rect 281062 38898 281146 39134
rect 281382 38898 281414 39134
rect 280794 3454 281414 38898
rect 280794 3218 280826 3454
rect 281062 3218 281146 3454
rect 281382 3218 281414 3454
rect 280794 3134 281414 3218
rect 280794 2898 280826 3134
rect 281062 2898 281146 3134
rect 281382 2898 281414 3134
rect 280794 -346 281414 2898
rect 280794 -582 280826 -346
rect 281062 -582 281146 -346
rect 281382 -582 281414 -346
rect 280794 -666 281414 -582
rect 280794 -902 280826 -666
rect 281062 -902 281146 -666
rect 281382 -902 281414 -666
rect 280794 -1894 281414 -902
rect 281954 680614 282574 711002
rect 291954 710598 292574 711590
rect 291954 710362 291986 710598
rect 292222 710362 292306 710598
rect 292542 710362 292574 710598
rect 291954 710278 292574 710362
rect 291954 710042 291986 710278
rect 292222 710042 292306 710278
rect 292542 710042 292574 710278
rect 288234 708678 288854 709670
rect 288234 708442 288266 708678
rect 288502 708442 288586 708678
rect 288822 708442 288854 708678
rect 288234 708358 288854 708442
rect 288234 708122 288266 708358
rect 288502 708122 288586 708358
rect 288822 708122 288854 708358
rect 281954 680378 281986 680614
rect 282222 680378 282306 680614
rect 282542 680378 282574 680614
rect 281954 680294 282574 680378
rect 281954 680058 281986 680294
rect 282222 680058 282306 680294
rect 282542 680058 282574 680294
rect 281954 644614 282574 680058
rect 281954 644378 281986 644614
rect 282222 644378 282306 644614
rect 282542 644378 282574 644614
rect 281954 644294 282574 644378
rect 281954 644058 281986 644294
rect 282222 644058 282306 644294
rect 282542 644058 282574 644294
rect 281954 608614 282574 644058
rect 281954 608378 281986 608614
rect 282222 608378 282306 608614
rect 282542 608378 282574 608614
rect 281954 608294 282574 608378
rect 281954 608058 281986 608294
rect 282222 608058 282306 608294
rect 282542 608058 282574 608294
rect 281954 572614 282574 608058
rect 281954 572378 281986 572614
rect 282222 572378 282306 572614
rect 282542 572378 282574 572614
rect 281954 572294 282574 572378
rect 281954 572058 281986 572294
rect 282222 572058 282306 572294
rect 282542 572058 282574 572294
rect 281954 536614 282574 572058
rect 281954 536378 281986 536614
rect 282222 536378 282306 536614
rect 282542 536378 282574 536614
rect 281954 536294 282574 536378
rect 281954 536058 281986 536294
rect 282222 536058 282306 536294
rect 282542 536058 282574 536294
rect 281954 500614 282574 536058
rect 281954 500378 281986 500614
rect 282222 500378 282306 500614
rect 282542 500378 282574 500614
rect 281954 500294 282574 500378
rect 281954 500058 281986 500294
rect 282222 500058 282306 500294
rect 282542 500058 282574 500294
rect 281954 464614 282574 500058
rect 281954 464378 281986 464614
rect 282222 464378 282306 464614
rect 282542 464378 282574 464614
rect 281954 464294 282574 464378
rect 281954 464058 281986 464294
rect 282222 464058 282306 464294
rect 282542 464058 282574 464294
rect 281954 428614 282574 464058
rect 281954 428378 281986 428614
rect 282222 428378 282306 428614
rect 282542 428378 282574 428614
rect 281954 428294 282574 428378
rect 281954 428058 281986 428294
rect 282222 428058 282306 428294
rect 282542 428058 282574 428294
rect 281954 392614 282574 428058
rect 281954 392378 281986 392614
rect 282222 392378 282306 392614
rect 282542 392378 282574 392614
rect 281954 392294 282574 392378
rect 281954 392058 281986 392294
rect 282222 392058 282306 392294
rect 282542 392058 282574 392294
rect 281954 356614 282574 392058
rect 281954 356378 281986 356614
rect 282222 356378 282306 356614
rect 282542 356378 282574 356614
rect 281954 356294 282574 356378
rect 281954 356058 281986 356294
rect 282222 356058 282306 356294
rect 282542 356058 282574 356294
rect 281954 320614 282574 356058
rect 281954 320378 281986 320614
rect 282222 320378 282306 320614
rect 282542 320378 282574 320614
rect 281954 320294 282574 320378
rect 281954 320058 281986 320294
rect 282222 320058 282306 320294
rect 282542 320058 282574 320294
rect 281954 284614 282574 320058
rect 281954 284378 281986 284614
rect 282222 284378 282306 284614
rect 282542 284378 282574 284614
rect 281954 284294 282574 284378
rect 281954 284058 281986 284294
rect 282222 284058 282306 284294
rect 282542 284058 282574 284294
rect 281954 248614 282574 284058
rect 281954 248378 281986 248614
rect 282222 248378 282306 248614
rect 282542 248378 282574 248614
rect 281954 248294 282574 248378
rect 281954 248058 281986 248294
rect 282222 248058 282306 248294
rect 282542 248058 282574 248294
rect 281954 212614 282574 248058
rect 281954 212378 281986 212614
rect 282222 212378 282306 212614
rect 282542 212378 282574 212614
rect 281954 212294 282574 212378
rect 281954 212058 281986 212294
rect 282222 212058 282306 212294
rect 282542 212058 282574 212294
rect 281954 176614 282574 212058
rect 281954 176378 281986 176614
rect 282222 176378 282306 176614
rect 282542 176378 282574 176614
rect 281954 176294 282574 176378
rect 281954 176058 281986 176294
rect 282222 176058 282306 176294
rect 282542 176058 282574 176294
rect 281954 140614 282574 176058
rect 281954 140378 281986 140614
rect 282222 140378 282306 140614
rect 282542 140378 282574 140614
rect 281954 140294 282574 140378
rect 281954 140058 281986 140294
rect 282222 140058 282306 140294
rect 282542 140058 282574 140294
rect 281954 104614 282574 140058
rect 281954 104378 281986 104614
rect 282222 104378 282306 104614
rect 282542 104378 282574 104614
rect 281954 104294 282574 104378
rect 281954 104058 281986 104294
rect 282222 104058 282306 104294
rect 282542 104058 282574 104294
rect 281954 68614 282574 104058
rect 281954 68378 281986 68614
rect 282222 68378 282306 68614
rect 282542 68378 282574 68614
rect 281954 68294 282574 68378
rect 281954 68058 281986 68294
rect 282222 68058 282306 68294
rect 282542 68058 282574 68294
rect 281954 32614 282574 68058
rect 281954 32378 281986 32614
rect 282222 32378 282306 32614
rect 282542 32378 282574 32614
rect 281954 32294 282574 32378
rect 281954 32058 281986 32294
rect 282222 32058 282306 32294
rect 282542 32058 282574 32294
rect 278234 -5382 278266 -5146
rect 278502 -5382 278586 -5146
rect 278822 -5382 278854 -5146
rect 278234 -5466 278854 -5382
rect 278234 -5702 278266 -5466
rect 278502 -5702 278586 -5466
rect 278822 -5702 278854 -5466
rect 278234 -5734 278854 -5702
rect 271954 -6342 271986 -6106
rect 272222 -6342 272306 -6106
rect 272542 -6342 272574 -6106
rect 271954 -6426 272574 -6342
rect 271954 -6662 271986 -6426
rect 272222 -6662 272306 -6426
rect 272542 -6662 272574 -6426
rect 271954 -7654 272574 -6662
rect 281954 -7066 282574 32058
rect 284514 706758 285134 707750
rect 284514 706522 284546 706758
rect 284782 706522 284866 706758
rect 285102 706522 285134 706758
rect 284514 706438 285134 706522
rect 284514 706202 284546 706438
rect 284782 706202 284866 706438
rect 285102 706202 285134 706438
rect 284514 691174 285134 706202
rect 284514 690938 284546 691174
rect 284782 690938 284866 691174
rect 285102 690938 285134 691174
rect 284514 690854 285134 690938
rect 284514 690618 284546 690854
rect 284782 690618 284866 690854
rect 285102 690618 285134 690854
rect 284514 655174 285134 690618
rect 284514 654938 284546 655174
rect 284782 654938 284866 655174
rect 285102 654938 285134 655174
rect 284514 654854 285134 654938
rect 284514 654618 284546 654854
rect 284782 654618 284866 654854
rect 285102 654618 285134 654854
rect 284514 619174 285134 654618
rect 284514 618938 284546 619174
rect 284782 618938 284866 619174
rect 285102 618938 285134 619174
rect 284514 618854 285134 618938
rect 284514 618618 284546 618854
rect 284782 618618 284866 618854
rect 285102 618618 285134 618854
rect 284514 583174 285134 618618
rect 284514 582938 284546 583174
rect 284782 582938 284866 583174
rect 285102 582938 285134 583174
rect 284514 582854 285134 582938
rect 284514 582618 284546 582854
rect 284782 582618 284866 582854
rect 285102 582618 285134 582854
rect 284514 547174 285134 582618
rect 284514 546938 284546 547174
rect 284782 546938 284866 547174
rect 285102 546938 285134 547174
rect 284514 546854 285134 546938
rect 284514 546618 284546 546854
rect 284782 546618 284866 546854
rect 285102 546618 285134 546854
rect 284514 511174 285134 546618
rect 284514 510938 284546 511174
rect 284782 510938 284866 511174
rect 285102 510938 285134 511174
rect 284514 510854 285134 510938
rect 284514 510618 284546 510854
rect 284782 510618 284866 510854
rect 285102 510618 285134 510854
rect 284514 475174 285134 510618
rect 284514 474938 284546 475174
rect 284782 474938 284866 475174
rect 285102 474938 285134 475174
rect 284514 474854 285134 474938
rect 284514 474618 284546 474854
rect 284782 474618 284866 474854
rect 285102 474618 285134 474854
rect 284514 439174 285134 474618
rect 284514 438938 284546 439174
rect 284782 438938 284866 439174
rect 285102 438938 285134 439174
rect 284514 438854 285134 438938
rect 284514 438618 284546 438854
rect 284782 438618 284866 438854
rect 285102 438618 285134 438854
rect 284514 403174 285134 438618
rect 284514 402938 284546 403174
rect 284782 402938 284866 403174
rect 285102 402938 285134 403174
rect 284514 402854 285134 402938
rect 284514 402618 284546 402854
rect 284782 402618 284866 402854
rect 285102 402618 285134 402854
rect 284514 367174 285134 402618
rect 284514 366938 284546 367174
rect 284782 366938 284866 367174
rect 285102 366938 285134 367174
rect 284514 366854 285134 366938
rect 284514 366618 284546 366854
rect 284782 366618 284866 366854
rect 285102 366618 285134 366854
rect 284514 331174 285134 366618
rect 284514 330938 284546 331174
rect 284782 330938 284866 331174
rect 285102 330938 285134 331174
rect 284514 330854 285134 330938
rect 284514 330618 284546 330854
rect 284782 330618 284866 330854
rect 285102 330618 285134 330854
rect 284514 295174 285134 330618
rect 284514 294938 284546 295174
rect 284782 294938 284866 295174
rect 285102 294938 285134 295174
rect 284514 294854 285134 294938
rect 284514 294618 284546 294854
rect 284782 294618 284866 294854
rect 285102 294618 285134 294854
rect 284514 259174 285134 294618
rect 284514 258938 284546 259174
rect 284782 258938 284866 259174
rect 285102 258938 285134 259174
rect 284514 258854 285134 258938
rect 284514 258618 284546 258854
rect 284782 258618 284866 258854
rect 285102 258618 285134 258854
rect 284514 223174 285134 258618
rect 284514 222938 284546 223174
rect 284782 222938 284866 223174
rect 285102 222938 285134 223174
rect 284514 222854 285134 222938
rect 284514 222618 284546 222854
rect 284782 222618 284866 222854
rect 285102 222618 285134 222854
rect 284514 187174 285134 222618
rect 284514 186938 284546 187174
rect 284782 186938 284866 187174
rect 285102 186938 285134 187174
rect 284514 186854 285134 186938
rect 284514 186618 284546 186854
rect 284782 186618 284866 186854
rect 285102 186618 285134 186854
rect 284514 151174 285134 186618
rect 284514 150938 284546 151174
rect 284782 150938 284866 151174
rect 285102 150938 285134 151174
rect 284514 150854 285134 150938
rect 284514 150618 284546 150854
rect 284782 150618 284866 150854
rect 285102 150618 285134 150854
rect 284514 115174 285134 150618
rect 284514 114938 284546 115174
rect 284782 114938 284866 115174
rect 285102 114938 285134 115174
rect 284514 114854 285134 114938
rect 284514 114618 284546 114854
rect 284782 114618 284866 114854
rect 285102 114618 285134 114854
rect 284514 79174 285134 114618
rect 284514 78938 284546 79174
rect 284782 78938 284866 79174
rect 285102 78938 285134 79174
rect 284514 78854 285134 78938
rect 284514 78618 284546 78854
rect 284782 78618 284866 78854
rect 285102 78618 285134 78854
rect 284514 43174 285134 78618
rect 284514 42938 284546 43174
rect 284782 42938 284866 43174
rect 285102 42938 285134 43174
rect 284514 42854 285134 42938
rect 284514 42618 284546 42854
rect 284782 42618 284866 42854
rect 285102 42618 285134 42854
rect 284514 7174 285134 42618
rect 284514 6938 284546 7174
rect 284782 6938 284866 7174
rect 285102 6938 285134 7174
rect 284514 6854 285134 6938
rect 284514 6618 284546 6854
rect 284782 6618 284866 6854
rect 285102 6618 285134 6854
rect 284514 -2266 285134 6618
rect 284514 -2502 284546 -2266
rect 284782 -2502 284866 -2266
rect 285102 -2502 285134 -2266
rect 284514 -2586 285134 -2502
rect 284514 -2822 284546 -2586
rect 284782 -2822 284866 -2586
rect 285102 -2822 285134 -2586
rect 284514 -3814 285134 -2822
rect 288234 694894 288854 708122
rect 288234 694658 288266 694894
rect 288502 694658 288586 694894
rect 288822 694658 288854 694894
rect 288234 694574 288854 694658
rect 288234 694338 288266 694574
rect 288502 694338 288586 694574
rect 288822 694338 288854 694574
rect 288234 658894 288854 694338
rect 288234 658658 288266 658894
rect 288502 658658 288586 658894
rect 288822 658658 288854 658894
rect 288234 658574 288854 658658
rect 288234 658338 288266 658574
rect 288502 658338 288586 658574
rect 288822 658338 288854 658574
rect 288234 622894 288854 658338
rect 288234 622658 288266 622894
rect 288502 622658 288586 622894
rect 288822 622658 288854 622894
rect 288234 622574 288854 622658
rect 288234 622338 288266 622574
rect 288502 622338 288586 622574
rect 288822 622338 288854 622574
rect 288234 586894 288854 622338
rect 288234 586658 288266 586894
rect 288502 586658 288586 586894
rect 288822 586658 288854 586894
rect 288234 586574 288854 586658
rect 288234 586338 288266 586574
rect 288502 586338 288586 586574
rect 288822 586338 288854 586574
rect 288234 550894 288854 586338
rect 288234 550658 288266 550894
rect 288502 550658 288586 550894
rect 288822 550658 288854 550894
rect 288234 550574 288854 550658
rect 288234 550338 288266 550574
rect 288502 550338 288586 550574
rect 288822 550338 288854 550574
rect 288234 514894 288854 550338
rect 288234 514658 288266 514894
rect 288502 514658 288586 514894
rect 288822 514658 288854 514894
rect 288234 514574 288854 514658
rect 288234 514338 288266 514574
rect 288502 514338 288586 514574
rect 288822 514338 288854 514574
rect 288234 478894 288854 514338
rect 288234 478658 288266 478894
rect 288502 478658 288586 478894
rect 288822 478658 288854 478894
rect 288234 478574 288854 478658
rect 288234 478338 288266 478574
rect 288502 478338 288586 478574
rect 288822 478338 288854 478574
rect 288234 442894 288854 478338
rect 288234 442658 288266 442894
rect 288502 442658 288586 442894
rect 288822 442658 288854 442894
rect 288234 442574 288854 442658
rect 288234 442338 288266 442574
rect 288502 442338 288586 442574
rect 288822 442338 288854 442574
rect 288234 406894 288854 442338
rect 288234 406658 288266 406894
rect 288502 406658 288586 406894
rect 288822 406658 288854 406894
rect 288234 406574 288854 406658
rect 288234 406338 288266 406574
rect 288502 406338 288586 406574
rect 288822 406338 288854 406574
rect 288234 370894 288854 406338
rect 288234 370658 288266 370894
rect 288502 370658 288586 370894
rect 288822 370658 288854 370894
rect 288234 370574 288854 370658
rect 288234 370338 288266 370574
rect 288502 370338 288586 370574
rect 288822 370338 288854 370574
rect 288234 334894 288854 370338
rect 288234 334658 288266 334894
rect 288502 334658 288586 334894
rect 288822 334658 288854 334894
rect 288234 334574 288854 334658
rect 288234 334338 288266 334574
rect 288502 334338 288586 334574
rect 288822 334338 288854 334574
rect 288234 298894 288854 334338
rect 288234 298658 288266 298894
rect 288502 298658 288586 298894
rect 288822 298658 288854 298894
rect 288234 298574 288854 298658
rect 288234 298338 288266 298574
rect 288502 298338 288586 298574
rect 288822 298338 288854 298574
rect 288234 262894 288854 298338
rect 288234 262658 288266 262894
rect 288502 262658 288586 262894
rect 288822 262658 288854 262894
rect 288234 262574 288854 262658
rect 288234 262338 288266 262574
rect 288502 262338 288586 262574
rect 288822 262338 288854 262574
rect 288234 226894 288854 262338
rect 288234 226658 288266 226894
rect 288502 226658 288586 226894
rect 288822 226658 288854 226894
rect 288234 226574 288854 226658
rect 288234 226338 288266 226574
rect 288502 226338 288586 226574
rect 288822 226338 288854 226574
rect 288234 190894 288854 226338
rect 288234 190658 288266 190894
rect 288502 190658 288586 190894
rect 288822 190658 288854 190894
rect 288234 190574 288854 190658
rect 288234 190338 288266 190574
rect 288502 190338 288586 190574
rect 288822 190338 288854 190574
rect 288234 154894 288854 190338
rect 288234 154658 288266 154894
rect 288502 154658 288586 154894
rect 288822 154658 288854 154894
rect 288234 154574 288854 154658
rect 288234 154338 288266 154574
rect 288502 154338 288586 154574
rect 288822 154338 288854 154574
rect 288234 118894 288854 154338
rect 288234 118658 288266 118894
rect 288502 118658 288586 118894
rect 288822 118658 288854 118894
rect 288234 118574 288854 118658
rect 288234 118338 288266 118574
rect 288502 118338 288586 118574
rect 288822 118338 288854 118574
rect 288234 82894 288854 118338
rect 288234 82658 288266 82894
rect 288502 82658 288586 82894
rect 288822 82658 288854 82894
rect 288234 82574 288854 82658
rect 288234 82338 288266 82574
rect 288502 82338 288586 82574
rect 288822 82338 288854 82574
rect 288234 46894 288854 82338
rect 288234 46658 288266 46894
rect 288502 46658 288586 46894
rect 288822 46658 288854 46894
rect 288234 46574 288854 46658
rect 288234 46338 288266 46574
rect 288502 46338 288586 46574
rect 288822 46338 288854 46574
rect 288234 10894 288854 46338
rect 288234 10658 288266 10894
rect 288502 10658 288586 10894
rect 288822 10658 288854 10894
rect 288234 10574 288854 10658
rect 288234 10338 288266 10574
rect 288502 10338 288586 10574
rect 288822 10338 288854 10574
rect 288234 -4186 288854 10338
rect 290794 705798 291414 705830
rect 290794 705562 290826 705798
rect 291062 705562 291146 705798
rect 291382 705562 291414 705798
rect 290794 705478 291414 705562
rect 290794 705242 290826 705478
rect 291062 705242 291146 705478
rect 291382 705242 291414 705478
rect 290794 669454 291414 705242
rect 290794 669218 290826 669454
rect 291062 669218 291146 669454
rect 291382 669218 291414 669454
rect 290794 669134 291414 669218
rect 290794 668898 290826 669134
rect 291062 668898 291146 669134
rect 291382 668898 291414 669134
rect 290794 633454 291414 668898
rect 290794 633218 290826 633454
rect 291062 633218 291146 633454
rect 291382 633218 291414 633454
rect 290794 633134 291414 633218
rect 290794 632898 290826 633134
rect 291062 632898 291146 633134
rect 291382 632898 291414 633134
rect 290794 597454 291414 632898
rect 290794 597218 290826 597454
rect 291062 597218 291146 597454
rect 291382 597218 291414 597454
rect 290794 597134 291414 597218
rect 290794 596898 290826 597134
rect 291062 596898 291146 597134
rect 291382 596898 291414 597134
rect 290794 561454 291414 596898
rect 290794 561218 290826 561454
rect 291062 561218 291146 561454
rect 291382 561218 291414 561454
rect 290794 561134 291414 561218
rect 290794 560898 290826 561134
rect 291062 560898 291146 561134
rect 291382 560898 291414 561134
rect 290794 525454 291414 560898
rect 290794 525218 290826 525454
rect 291062 525218 291146 525454
rect 291382 525218 291414 525454
rect 290794 525134 291414 525218
rect 290794 524898 290826 525134
rect 291062 524898 291146 525134
rect 291382 524898 291414 525134
rect 290794 489454 291414 524898
rect 290794 489218 290826 489454
rect 291062 489218 291146 489454
rect 291382 489218 291414 489454
rect 290794 489134 291414 489218
rect 290794 488898 290826 489134
rect 291062 488898 291146 489134
rect 291382 488898 291414 489134
rect 290794 453454 291414 488898
rect 290794 453218 290826 453454
rect 291062 453218 291146 453454
rect 291382 453218 291414 453454
rect 290794 453134 291414 453218
rect 290794 452898 290826 453134
rect 291062 452898 291146 453134
rect 291382 452898 291414 453134
rect 290794 417454 291414 452898
rect 290794 417218 290826 417454
rect 291062 417218 291146 417454
rect 291382 417218 291414 417454
rect 290794 417134 291414 417218
rect 290794 416898 290826 417134
rect 291062 416898 291146 417134
rect 291382 416898 291414 417134
rect 290794 381454 291414 416898
rect 290794 381218 290826 381454
rect 291062 381218 291146 381454
rect 291382 381218 291414 381454
rect 290794 381134 291414 381218
rect 290794 380898 290826 381134
rect 291062 380898 291146 381134
rect 291382 380898 291414 381134
rect 290794 345454 291414 380898
rect 290794 345218 290826 345454
rect 291062 345218 291146 345454
rect 291382 345218 291414 345454
rect 290794 345134 291414 345218
rect 290794 344898 290826 345134
rect 291062 344898 291146 345134
rect 291382 344898 291414 345134
rect 290794 309454 291414 344898
rect 290794 309218 290826 309454
rect 291062 309218 291146 309454
rect 291382 309218 291414 309454
rect 290794 309134 291414 309218
rect 290794 308898 290826 309134
rect 291062 308898 291146 309134
rect 291382 308898 291414 309134
rect 290794 273454 291414 308898
rect 290794 273218 290826 273454
rect 291062 273218 291146 273454
rect 291382 273218 291414 273454
rect 290794 273134 291414 273218
rect 290794 272898 290826 273134
rect 291062 272898 291146 273134
rect 291382 272898 291414 273134
rect 290794 237454 291414 272898
rect 290794 237218 290826 237454
rect 291062 237218 291146 237454
rect 291382 237218 291414 237454
rect 290794 237134 291414 237218
rect 290794 236898 290826 237134
rect 291062 236898 291146 237134
rect 291382 236898 291414 237134
rect 290794 201454 291414 236898
rect 290794 201218 290826 201454
rect 291062 201218 291146 201454
rect 291382 201218 291414 201454
rect 290794 201134 291414 201218
rect 290794 200898 290826 201134
rect 291062 200898 291146 201134
rect 291382 200898 291414 201134
rect 290794 165454 291414 200898
rect 290794 165218 290826 165454
rect 291062 165218 291146 165454
rect 291382 165218 291414 165454
rect 290794 165134 291414 165218
rect 290794 164898 290826 165134
rect 291062 164898 291146 165134
rect 291382 164898 291414 165134
rect 290794 129454 291414 164898
rect 290794 129218 290826 129454
rect 291062 129218 291146 129454
rect 291382 129218 291414 129454
rect 290794 129134 291414 129218
rect 290794 128898 290826 129134
rect 291062 128898 291146 129134
rect 291382 128898 291414 129134
rect 290794 93454 291414 128898
rect 290794 93218 290826 93454
rect 291062 93218 291146 93454
rect 291382 93218 291414 93454
rect 290794 93134 291414 93218
rect 290794 92898 290826 93134
rect 291062 92898 291146 93134
rect 291382 92898 291414 93134
rect 290794 57454 291414 92898
rect 290794 57218 290826 57454
rect 291062 57218 291146 57454
rect 291382 57218 291414 57454
rect 290794 57134 291414 57218
rect 290794 56898 290826 57134
rect 291062 56898 291146 57134
rect 291382 56898 291414 57134
rect 290794 21454 291414 56898
rect 290794 21218 290826 21454
rect 291062 21218 291146 21454
rect 291382 21218 291414 21454
rect 290794 21134 291414 21218
rect 290794 20898 290826 21134
rect 291062 20898 291146 21134
rect 291382 20898 291414 21134
rect 290794 -1306 291414 20898
rect 290794 -1542 290826 -1306
rect 291062 -1542 291146 -1306
rect 291382 -1542 291414 -1306
rect 290794 -1626 291414 -1542
rect 290794 -1862 290826 -1626
rect 291062 -1862 291146 -1626
rect 291382 -1862 291414 -1626
rect 290794 -1894 291414 -1862
rect 291954 698614 292574 710042
rect 301954 711558 302574 711590
rect 301954 711322 301986 711558
rect 302222 711322 302306 711558
rect 302542 711322 302574 711558
rect 301954 711238 302574 711322
rect 301954 711002 301986 711238
rect 302222 711002 302306 711238
rect 302542 711002 302574 711238
rect 298234 709638 298854 709670
rect 298234 709402 298266 709638
rect 298502 709402 298586 709638
rect 298822 709402 298854 709638
rect 298234 709318 298854 709402
rect 298234 709082 298266 709318
rect 298502 709082 298586 709318
rect 298822 709082 298854 709318
rect 291954 698378 291986 698614
rect 292222 698378 292306 698614
rect 292542 698378 292574 698614
rect 291954 698294 292574 698378
rect 291954 698058 291986 698294
rect 292222 698058 292306 698294
rect 292542 698058 292574 698294
rect 291954 662614 292574 698058
rect 291954 662378 291986 662614
rect 292222 662378 292306 662614
rect 292542 662378 292574 662614
rect 291954 662294 292574 662378
rect 291954 662058 291986 662294
rect 292222 662058 292306 662294
rect 292542 662058 292574 662294
rect 291954 626614 292574 662058
rect 291954 626378 291986 626614
rect 292222 626378 292306 626614
rect 292542 626378 292574 626614
rect 291954 626294 292574 626378
rect 291954 626058 291986 626294
rect 292222 626058 292306 626294
rect 292542 626058 292574 626294
rect 291954 590614 292574 626058
rect 291954 590378 291986 590614
rect 292222 590378 292306 590614
rect 292542 590378 292574 590614
rect 291954 590294 292574 590378
rect 291954 590058 291986 590294
rect 292222 590058 292306 590294
rect 292542 590058 292574 590294
rect 291954 554614 292574 590058
rect 291954 554378 291986 554614
rect 292222 554378 292306 554614
rect 292542 554378 292574 554614
rect 291954 554294 292574 554378
rect 291954 554058 291986 554294
rect 292222 554058 292306 554294
rect 292542 554058 292574 554294
rect 291954 518614 292574 554058
rect 291954 518378 291986 518614
rect 292222 518378 292306 518614
rect 292542 518378 292574 518614
rect 291954 518294 292574 518378
rect 291954 518058 291986 518294
rect 292222 518058 292306 518294
rect 292542 518058 292574 518294
rect 291954 482614 292574 518058
rect 291954 482378 291986 482614
rect 292222 482378 292306 482614
rect 292542 482378 292574 482614
rect 291954 482294 292574 482378
rect 291954 482058 291986 482294
rect 292222 482058 292306 482294
rect 292542 482058 292574 482294
rect 291954 446614 292574 482058
rect 291954 446378 291986 446614
rect 292222 446378 292306 446614
rect 292542 446378 292574 446614
rect 291954 446294 292574 446378
rect 291954 446058 291986 446294
rect 292222 446058 292306 446294
rect 292542 446058 292574 446294
rect 291954 410614 292574 446058
rect 291954 410378 291986 410614
rect 292222 410378 292306 410614
rect 292542 410378 292574 410614
rect 291954 410294 292574 410378
rect 291954 410058 291986 410294
rect 292222 410058 292306 410294
rect 292542 410058 292574 410294
rect 291954 374614 292574 410058
rect 291954 374378 291986 374614
rect 292222 374378 292306 374614
rect 292542 374378 292574 374614
rect 291954 374294 292574 374378
rect 291954 374058 291986 374294
rect 292222 374058 292306 374294
rect 292542 374058 292574 374294
rect 291954 338614 292574 374058
rect 291954 338378 291986 338614
rect 292222 338378 292306 338614
rect 292542 338378 292574 338614
rect 291954 338294 292574 338378
rect 291954 338058 291986 338294
rect 292222 338058 292306 338294
rect 292542 338058 292574 338294
rect 291954 302614 292574 338058
rect 291954 302378 291986 302614
rect 292222 302378 292306 302614
rect 292542 302378 292574 302614
rect 291954 302294 292574 302378
rect 291954 302058 291986 302294
rect 292222 302058 292306 302294
rect 292542 302058 292574 302294
rect 291954 266614 292574 302058
rect 291954 266378 291986 266614
rect 292222 266378 292306 266614
rect 292542 266378 292574 266614
rect 291954 266294 292574 266378
rect 291954 266058 291986 266294
rect 292222 266058 292306 266294
rect 292542 266058 292574 266294
rect 291954 230614 292574 266058
rect 291954 230378 291986 230614
rect 292222 230378 292306 230614
rect 292542 230378 292574 230614
rect 291954 230294 292574 230378
rect 291954 230058 291986 230294
rect 292222 230058 292306 230294
rect 292542 230058 292574 230294
rect 291954 194614 292574 230058
rect 291954 194378 291986 194614
rect 292222 194378 292306 194614
rect 292542 194378 292574 194614
rect 291954 194294 292574 194378
rect 291954 194058 291986 194294
rect 292222 194058 292306 194294
rect 292542 194058 292574 194294
rect 291954 158614 292574 194058
rect 291954 158378 291986 158614
rect 292222 158378 292306 158614
rect 292542 158378 292574 158614
rect 291954 158294 292574 158378
rect 291954 158058 291986 158294
rect 292222 158058 292306 158294
rect 292542 158058 292574 158294
rect 291954 122614 292574 158058
rect 291954 122378 291986 122614
rect 292222 122378 292306 122614
rect 292542 122378 292574 122614
rect 291954 122294 292574 122378
rect 291954 122058 291986 122294
rect 292222 122058 292306 122294
rect 292542 122058 292574 122294
rect 291954 86614 292574 122058
rect 291954 86378 291986 86614
rect 292222 86378 292306 86614
rect 292542 86378 292574 86614
rect 291954 86294 292574 86378
rect 291954 86058 291986 86294
rect 292222 86058 292306 86294
rect 292542 86058 292574 86294
rect 291954 50614 292574 86058
rect 291954 50378 291986 50614
rect 292222 50378 292306 50614
rect 292542 50378 292574 50614
rect 291954 50294 292574 50378
rect 291954 50058 291986 50294
rect 292222 50058 292306 50294
rect 292542 50058 292574 50294
rect 291954 14614 292574 50058
rect 291954 14378 291986 14614
rect 292222 14378 292306 14614
rect 292542 14378 292574 14614
rect 291954 14294 292574 14378
rect 291954 14058 291986 14294
rect 292222 14058 292306 14294
rect 292542 14058 292574 14294
rect 288234 -4422 288266 -4186
rect 288502 -4422 288586 -4186
rect 288822 -4422 288854 -4186
rect 288234 -4506 288854 -4422
rect 288234 -4742 288266 -4506
rect 288502 -4742 288586 -4506
rect 288822 -4742 288854 -4506
rect 288234 -5734 288854 -4742
rect 281954 -7302 281986 -7066
rect 282222 -7302 282306 -7066
rect 282542 -7302 282574 -7066
rect 281954 -7386 282574 -7302
rect 281954 -7622 281986 -7386
rect 282222 -7622 282306 -7386
rect 282542 -7622 282574 -7386
rect 281954 -7654 282574 -7622
rect 291954 -6106 292574 14058
rect 294514 707718 295134 707750
rect 294514 707482 294546 707718
rect 294782 707482 294866 707718
rect 295102 707482 295134 707718
rect 294514 707398 295134 707482
rect 294514 707162 294546 707398
rect 294782 707162 294866 707398
rect 295102 707162 295134 707398
rect 294514 673174 295134 707162
rect 294514 672938 294546 673174
rect 294782 672938 294866 673174
rect 295102 672938 295134 673174
rect 294514 672854 295134 672938
rect 294514 672618 294546 672854
rect 294782 672618 294866 672854
rect 295102 672618 295134 672854
rect 294514 637174 295134 672618
rect 294514 636938 294546 637174
rect 294782 636938 294866 637174
rect 295102 636938 295134 637174
rect 294514 636854 295134 636938
rect 294514 636618 294546 636854
rect 294782 636618 294866 636854
rect 295102 636618 295134 636854
rect 294514 601174 295134 636618
rect 294514 600938 294546 601174
rect 294782 600938 294866 601174
rect 295102 600938 295134 601174
rect 294514 600854 295134 600938
rect 294514 600618 294546 600854
rect 294782 600618 294866 600854
rect 295102 600618 295134 600854
rect 294514 565174 295134 600618
rect 294514 564938 294546 565174
rect 294782 564938 294866 565174
rect 295102 564938 295134 565174
rect 294514 564854 295134 564938
rect 294514 564618 294546 564854
rect 294782 564618 294866 564854
rect 295102 564618 295134 564854
rect 294514 529174 295134 564618
rect 294514 528938 294546 529174
rect 294782 528938 294866 529174
rect 295102 528938 295134 529174
rect 294514 528854 295134 528938
rect 294514 528618 294546 528854
rect 294782 528618 294866 528854
rect 295102 528618 295134 528854
rect 294514 493174 295134 528618
rect 294514 492938 294546 493174
rect 294782 492938 294866 493174
rect 295102 492938 295134 493174
rect 294514 492854 295134 492938
rect 294514 492618 294546 492854
rect 294782 492618 294866 492854
rect 295102 492618 295134 492854
rect 294514 457174 295134 492618
rect 294514 456938 294546 457174
rect 294782 456938 294866 457174
rect 295102 456938 295134 457174
rect 294514 456854 295134 456938
rect 294514 456618 294546 456854
rect 294782 456618 294866 456854
rect 295102 456618 295134 456854
rect 294514 421174 295134 456618
rect 294514 420938 294546 421174
rect 294782 420938 294866 421174
rect 295102 420938 295134 421174
rect 294514 420854 295134 420938
rect 294514 420618 294546 420854
rect 294782 420618 294866 420854
rect 295102 420618 295134 420854
rect 294514 385174 295134 420618
rect 294514 384938 294546 385174
rect 294782 384938 294866 385174
rect 295102 384938 295134 385174
rect 294514 384854 295134 384938
rect 294514 384618 294546 384854
rect 294782 384618 294866 384854
rect 295102 384618 295134 384854
rect 294514 349174 295134 384618
rect 294514 348938 294546 349174
rect 294782 348938 294866 349174
rect 295102 348938 295134 349174
rect 294514 348854 295134 348938
rect 294514 348618 294546 348854
rect 294782 348618 294866 348854
rect 295102 348618 295134 348854
rect 294514 313174 295134 348618
rect 294514 312938 294546 313174
rect 294782 312938 294866 313174
rect 295102 312938 295134 313174
rect 294514 312854 295134 312938
rect 294514 312618 294546 312854
rect 294782 312618 294866 312854
rect 295102 312618 295134 312854
rect 294514 277174 295134 312618
rect 294514 276938 294546 277174
rect 294782 276938 294866 277174
rect 295102 276938 295134 277174
rect 294514 276854 295134 276938
rect 294514 276618 294546 276854
rect 294782 276618 294866 276854
rect 295102 276618 295134 276854
rect 294514 241174 295134 276618
rect 294514 240938 294546 241174
rect 294782 240938 294866 241174
rect 295102 240938 295134 241174
rect 294514 240854 295134 240938
rect 294514 240618 294546 240854
rect 294782 240618 294866 240854
rect 295102 240618 295134 240854
rect 294514 205174 295134 240618
rect 294514 204938 294546 205174
rect 294782 204938 294866 205174
rect 295102 204938 295134 205174
rect 294514 204854 295134 204938
rect 294514 204618 294546 204854
rect 294782 204618 294866 204854
rect 295102 204618 295134 204854
rect 294514 169174 295134 204618
rect 294514 168938 294546 169174
rect 294782 168938 294866 169174
rect 295102 168938 295134 169174
rect 294514 168854 295134 168938
rect 294514 168618 294546 168854
rect 294782 168618 294866 168854
rect 295102 168618 295134 168854
rect 294514 133174 295134 168618
rect 294514 132938 294546 133174
rect 294782 132938 294866 133174
rect 295102 132938 295134 133174
rect 294514 132854 295134 132938
rect 294514 132618 294546 132854
rect 294782 132618 294866 132854
rect 295102 132618 295134 132854
rect 294514 97174 295134 132618
rect 294514 96938 294546 97174
rect 294782 96938 294866 97174
rect 295102 96938 295134 97174
rect 294514 96854 295134 96938
rect 294514 96618 294546 96854
rect 294782 96618 294866 96854
rect 295102 96618 295134 96854
rect 294514 61174 295134 96618
rect 294514 60938 294546 61174
rect 294782 60938 294866 61174
rect 295102 60938 295134 61174
rect 294514 60854 295134 60938
rect 294514 60618 294546 60854
rect 294782 60618 294866 60854
rect 295102 60618 295134 60854
rect 294514 25174 295134 60618
rect 294514 24938 294546 25174
rect 294782 24938 294866 25174
rect 295102 24938 295134 25174
rect 294514 24854 295134 24938
rect 294514 24618 294546 24854
rect 294782 24618 294866 24854
rect 295102 24618 295134 24854
rect 294514 -3226 295134 24618
rect 294514 -3462 294546 -3226
rect 294782 -3462 294866 -3226
rect 295102 -3462 295134 -3226
rect 294514 -3546 295134 -3462
rect 294514 -3782 294546 -3546
rect 294782 -3782 294866 -3546
rect 295102 -3782 295134 -3546
rect 294514 -3814 295134 -3782
rect 298234 676894 298854 709082
rect 298234 676658 298266 676894
rect 298502 676658 298586 676894
rect 298822 676658 298854 676894
rect 298234 676574 298854 676658
rect 298234 676338 298266 676574
rect 298502 676338 298586 676574
rect 298822 676338 298854 676574
rect 298234 640894 298854 676338
rect 298234 640658 298266 640894
rect 298502 640658 298586 640894
rect 298822 640658 298854 640894
rect 298234 640574 298854 640658
rect 298234 640338 298266 640574
rect 298502 640338 298586 640574
rect 298822 640338 298854 640574
rect 298234 604894 298854 640338
rect 298234 604658 298266 604894
rect 298502 604658 298586 604894
rect 298822 604658 298854 604894
rect 298234 604574 298854 604658
rect 298234 604338 298266 604574
rect 298502 604338 298586 604574
rect 298822 604338 298854 604574
rect 298234 568894 298854 604338
rect 298234 568658 298266 568894
rect 298502 568658 298586 568894
rect 298822 568658 298854 568894
rect 298234 568574 298854 568658
rect 298234 568338 298266 568574
rect 298502 568338 298586 568574
rect 298822 568338 298854 568574
rect 298234 532894 298854 568338
rect 298234 532658 298266 532894
rect 298502 532658 298586 532894
rect 298822 532658 298854 532894
rect 298234 532574 298854 532658
rect 298234 532338 298266 532574
rect 298502 532338 298586 532574
rect 298822 532338 298854 532574
rect 298234 496894 298854 532338
rect 298234 496658 298266 496894
rect 298502 496658 298586 496894
rect 298822 496658 298854 496894
rect 298234 496574 298854 496658
rect 298234 496338 298266 496574
rect 298502 496338 298586 496574
rect 298822 496338 298854 496574
rect 298234 460894 298854 496338
rect 298234 460658 298266 460894
rect 298502 460658 298586 460894
rect 298822 460658 298854 460894
rect 298234 460574 298854 460658
rect 298234 460338 298266 460574
rect 298502 460338 298586 460574
rect 298822 460338 298854 460574
rect 298234 424894 298854 460338
rect 298234 424658 298266 424894
rect 298502 424658 298586 424894
rect 298822 424658 298854 424894
rect 298234 424574 298854 424658
rect 298234 424338 298266 424574
rect 298502 424338 298586 424574
rect 298822 424338 298854 424574
rect 298234 388894 298854 424338
rect 298234 388658 298266 388894
rect 298502 388658 298586 388894
rect 298822 388658 298854 388894
rect 298234 388574 298854 388658
rect 298234 388338 298266 388574
rect 298502 388338 298586 388574
rect 298822 388338 298854 388574
rect 298234 352894 298854 388338
rect 298234 352658 298266 352894
rect 298502 352658 298586 352894
rect 298822 352658 298854 352894
rect 298234 352574 298854 352658
rect 298234 352338 298266 352574
rect 298502 352338 298586 352574
rect 298822 352338 298854 352574
rect 298234 316894 298854 352338
rect 298234 316658 298266 316894
rect 298502 316658 298586 316894
rect 298822 316658 298854 316894
rect 298234 316574 298854 316658
rect 298234 316338 298266 316574
rect 298502 316338 298586 316574
rect 298822 316338 298854 316574
rect 298234 280894 298854 316338
rect 298234 280658 298266 280894
rect 298502 280658 298586 280894
rect 298822 280658 298854 280894
rect 298234 280574 298854 280658
rect 298234 280338 298266 280574
rect 298502 280338 298586 280574
rect 298822 280338 298854 280574
rect 298234 244894 298854 280338
rect 298234 244658 298266 244894
rect 298502 244658 298586 244894
rect 298822 244658 298854 244894
rect 298234 244574 298854 244658
rect 298234 244338 298266 244574
rect 298502 244338 298586 244574
rect 298822 244338 298854 244574
rect 298234 208894 298854 244338
rect 298234 208658 298266 208894
rect 298502 208658 298586 208894
rect 298822 208658 298854 208894
rect 298234 208574 298854 208658
rect 298234 208338 298266 208574
rect 298502 208338 298586 208574
rect 298822 208338 298854 208574
rect 298234 172894 298854 208338
rect 298234 172658 298266 172894
rect 298502 172658 298586 172894
rect 298822 172658 298854 172894
rect 298234 172574 298854 172658
rect 298234 172338 298266 172574
rect 298502 172338 298586 172574
rect 298822 172338 298854 172574
rect 298234 136894 298854 172338
rect 298234 136658 298266 136894
rect 298502 136658 298586 136894
rect 298822 136658 298854 136894
rect 298234 136574 298854 136658
rect 298234 136338 298266 136574
rect 298502 136338 298586 136574
rect 298822 136338 298854 136574
rect 298234 100894 298854 136338
rect 298234 100658 298266 100894
rect 298502 100658 298586 100894
rect 298822 100658 298854 100894
rect 298234 100574 298854 100658
rect 298234 100338 298266 100574
rect 298502 100338 298586 100574
rect 298822 100338 298854 100574
rect 298234 64894 298854 100338
rect 298234 64658 298266 64894
rect 298502 64658 298586 64894
rect 298822 64658 298854 64894
rect 298234 64574 298854 64658
rect 298234 64338 298266 64574
rect 298502 64338 298586 64574
rect 298822 64338 298854 64574
rect 298234 28894 298854 64338
rect 298234 28658 298266 28894
rect 298502 28658 298586 28894
rect 298822 28658 298854 28894
rect 298234 28574 298854 28658
rect 298234 28338 298266 28574
rect 298502 28338 298586 28574
rect 298822 28338 298854 28574
rect 298234 -5146 298854 28338
rect 300794 704838 301414 705830
rect 300794 704602 300826 704838
rect 301062 704602 301146 704838
rect 301382 704602 301414 704838
rect 300794 704518 301414 704602
rect 300794 704282 300826 704518
rect 301062 704282 301146 704518
rect 301382 704282 301414 704518
rect 300794 687454 301414 704282
rect 300794 687218 300826 687454
rect 301062 687218 301146 687454
rect 301382 687218 301414 687454
rect 300794 687134 301414 687218
rect 300794 686898 300826 687134
rect 301062 686898 301146 687134
rect 301382 686898 301414 687134
rect 300794 651454 301414 686898
rect 300794 651218 300826 651454
rect 301062 651218 301146 651454
rect 301382 651218 301414 651454
rect 300794 651134 301414 651218
rect 300794 650898 300826 651134
rect 301062 650898 301146 651134
rect 301382 650898 301414 651134
rect 300794 615454 301414 650898
rect 300794 615218 300826 615454
rect 301062 615218 301146 615454
rect 301382 615218 301414 615454
rect 300794 615134 301414 615218
rect 300794 614898 300826 615134
rect 301062 614898 301146 615134
rect 301382 614898 301414 615134
rect 300794 579454 301414 614898
rect 300794 579218 300826 579454
rect 301062 579218 301146 579454
rect 301382 579218 301414 579454
rect 300794 579134 301414 579218
rect 300794 578898 300826 579134
rect 301062 578898 301146 579134
rect 301382 578898 301414 579134
rect 300794 543454 301414 578898
rect 300794 543218 300826 543454
rect 301062 543218 301146 543454
rect 301382 543218 301414 543454
rect 300794 543134 301414 543218
rect 300794 542898 300826 543134
rect 301062 542898 301146 543134
rect 301382 542898 301414 543134
rect 300794 507454 301414 542898
rect 300794 507218 300826 507454
rect 301062 507218 301146 507454
rect 301382 507218 301414 507454
rect 300794 507134 301414 507218
rect 300794 506898 300826 507134
rect 301062 506898 301146 507134
rect 301382 506898 301414 507134
rect 300794 471454 301414 506898
rect 300794 471218 300826 471454
rect 301062 471218 301146 471454
rect 301382 471218 301414 471454
rect 300794 471134 301414 471218
rect 300794 470898 300826 471134
rect 301062 470898 301146 471134
rect 301382 470898 301414 471134
rect 300794 435454 301414 470898
rect 300794 435218 300826 435454
rect 301062 435218 301146 435454
rect 301382 435218 301414 435454
rect 300794 435134 301414 435218
rect 300794 434898 300826 435134
rect 301062 434898 301146 435134
rect 301382 434898 301414 435134
rect 300794 399454 301414 434898
rect 300794 399218 300826 399454
rect 301062 399218 301146 399454
rect 301382 399218 301414 399454
rect 300794 399134 301414 399218
rect 300794 398898 300826 399134
rect 301062 398898 301146 399134
rect 301382 398898 301414 399134
rect 300794 363454 301414 398898
rect 300794 363218 300826 363454
rect 301062 363218 301146 363454
rect 301382 363218 301414 363454
rect 300794 363134 301414 363218
rect 300794 362898 300826 363134
rect 301062 362898 301146 363134
rect 301382 362898 301414 363134
rect 300794 327454 301414 362898
rect 300794 327218 300826 327454
rect 301062 327218 301146 327454
rect 301382 327218 301414 327454
rect 300794 327134 301414 327218
rect 300794 326898 300826 327134
rect 301062 326898 301146 327134
rect 301382 326898 301414 327134
rect 300794 291454 301414 326898
rect 300794 291218 300826 291454
rect 301062 291218 301146 291454
rect 301382 291218 301414 291454
rect 300794 291134 301414 291218
rect 300794 290898 300826 291134
rect 301062 290898 301146 291134
rect 301382 290898 301414 291134
rect 300794 255454 301414 290898
rect 300794 255218 300826 255454
rect 301062 255218 301146 255454
rect 301382 255218 301414 255454
rect 300794 255134 301414 255218
rect 300794 254898 300826 255134
rect 301062 254898 301146 255134
rect 301382 254898 301414 255134
rect 300794 219454 301414 254898
rect 300794 219218 300826 219454
rect 301062 219218 301146 219454
rect 301382 219218 301414 219454
rect 300794 219134 301414 219218
rect 300794 218898 300826 219134
rect 301062 218898 301146 219134
rect 301382 218898 301414 219134
rect 300794 183454 301414 218898
rect 300794 183218 300826 183454
rect 301062 183218 301146 183454
rect 301382 183218 301414 183454
rect 300794 183134 301414 183218
rect 300794 182898 300826 183134
rect 301062 182898 301146 183134
rect 301382 182898 301414 183134
rect 300794 147454 301414 182898
rect 300794 147218 300826 147454
rect 301062 147218 301146 147454
rect 301382 147218 301414 147454
rect 300794 147134 301414 147218
rect 300794 146898 300826 147134
rect 301062 146898 301146 147134
rect 301382 146898 301414 147134
rect 300794 111454 301414 146898
rect 300794 111218 300826 111454
rect 301062 111218 301146 111454
rect 301382 111218 301414 111454
rect 300794 111134 301414 111218
rect 300794 110898 300826 111134
rect 301062 110898 301146 111134
rect 301382 110898 301414 111134
rect 300794 75454 301414 110898
rect 300794 75218 300826 75454
rect 301062 75218 301146 75454
rect 301382 75218 301414 75454
rect 300794 75134 301414 75218
rect 300794 74898 300826 75134
rect 301062 74898 301146 75134
rect 301382 74898 301414 75134
rect 300794 39454 301414 74898
rect 300794 39218 300826 39454
rect 301062 39218 301146 39454
rect 301382 39218 301414 39454
rect 300794 39134 301414 39218
rect 300794 38898 300826 39134
rect 301062 38898 301146 39134
rect 301382 38898 301414 39134
rect 300794 3454 301414 38898
rect 300794 3218 300826 3454
rect 301062 3218 301146 3454
rect 301382 3218 301414 3454
rect 300794 3134 301414 3218
rect 300794 2898 300826 3134
rect 301062 2898 301146 3134
rect 301382 2898 301414 3134
rect 300794 -346 301414 2898
rect 300794 -582 300826 -346
rect 301062 -582 301146 -346
rect 301382 -582 301414 -346
rect 300794 -666 301414 -582
rect 300794 -902 300826 -666
rect 301062 -902 301146 -666
rect 301382 -902 301414 -666
rect 300794 -1894 301414 -902
rect 301954 680614 302574 711002
rect 311954 710598 312574 711590
rect 311954 710362 311986 710598
rect 312222 710362 312306 710598
rect 312542 710362 312574 710598
rect 311954 710278 312574 710362
rect 311954 710042 311986 710278
rect 312222 710042 312306 710278
rect 312542 710042 312574 710278
rect 308234 708678 308854 709670
rect 308234 708442 308266 708678
rect 308502 708442 308586 708678
rect 308822 708442 308854 708678
rect 308234 708358 308854 708442
rect 308234 708122 308266 708358
rect 308502 708122 308586 708358
rect 308822 708122 308854 708358
rect 301954 680378 301986 680614
rect 302222 680378 302306 680614
rect 302542 680378 302574 680614
rect 301954 680294 302574 680378
rect 301954 680058 301986 680294
rect 302222 680058 302306 680294
rect 302542 680058 302574 680294
rect 301954 644614 302574 680058
rect 301954 644378 301986 644614
rect 302222 644378 302306 644614
rect 302542 644378 302574 644614
rect 301954 644294 302574 644378
rect 301954 644058 301986 644294
rect 302222 644058 302306 644294
rect 302542 644058 302574 644294
rect 301954 608614 302574 644058
rect 301954 608378 301986 608614
rect 302222 608378 302306 608614
rect 302542 608378 302574 608614
rect 301954 608294 302574 608378
rect 301954 608058 301986 608294
rect 302222 608058 302306 608294
rect 302542 608058 302574 608294
rect 301954 572614 302574 608058
rect 301954 572378 301986 572614
rect 302222 572378 302306 572614
rect 302542 572378 302574 572614
rect 301954 572294 302574 572378
rect 301954 572058 301986 572294
rect 302222 572058 302306 572294
rect 302542 572058 302574 572294
rect 301954 536614 302574 572058
rect 301954 536378 301986 536614
rect 302222 536378 302306 536614
rect 302542 536378 302574 536614
rect 301954 536294 302574 536378
rect 301954 536058 301986 536294
rect 302222 536058 302306 536294
rect 302542 536058 302574 536294
rect 301954 500614 302574 536058
rect 301954 500378 301986 500614
rect 302222 500378 302306 500614
rect 302542 500378 302574 500614
rect 301954 500294 302574 500378
rect 301954 500058 301986 500294
rect 302222 500058 302306 500294
rect 302542 500058 302574 500294
rect 301954 464614 302574 500058
rect 301954 464378 301986 464614
rect 302222 464378 302306 464614
rect 302542 464378 302574 464614
rect 301954 464294 302574 464378
rect 301954 464058 301986 464294
rect 302222 464058 302306 464294
rect 302542 464058 302574 464294
rect 301954 428614 302574 464058
rect 301954 428378 301986 428614
rect 302222 428378 302306 428614
rect 302542 428378 302574 428614
rect 301954 428294 302574 428378
rect 301954 428058 301986 428294
rect 302222 428058 302306 428294
rect 302542 428058 302574 428294
rect 301954 392614 302574 428058
rect 301954 392378 301986 392614
rect 302222 392378 302306 392614
rect 302542 392378 302574 392614
rect 301954 392294 302574 392378
rect 301954 392058 301986 392294
rect 302222 392058 302306 392294
rect 302542 392058 302574 392294
rect 301954 356614 302574 392058
rect 301954 356378 301986 356614
rect 302222 356378 302306 356614
rect 302542 356378 302574 356614
rect 301954 356294 302574 356378
rect 301954 356058 301986 356294
rect 302222 356058 302306 356294
rect 302542 356058 302574 356294
rect 301954 320614 302574 356058
rect 301954 320378 301986 320614
rect 302222 320378 302306 320614
rect 302542 320378 302574 320614
rect 301954 320294 302574 320378
rect 301954 320058 301986 320294
rect 302222 320058 302306 320294
rect 302542 320058 302574 320294
rect 301954 284614 302574 320058
rect 301954 284378 301986 284614
rect 302222 284378 302306 284614
rect 302542 284378 302574 284614
rect 301954 284294 302574 284378
rect 301954 284058 301986 284294
rect 302222 284058 302306 284294
rect 302542 284058 302574 284294
rect 301954 248614 302574 284058
rect 301954 248378 301986 248614
rect 302222 248378 302306 248614
rect 302542 248378 302574 248614
rect 301954 248294 302574 248378
rect 301954 248058 301986 248294
rect 302222 248058 302306 248294
rect 302542 248058 302574 248294
rect 301954 212614 302574 248058
rect 301954 212378 301986 212614
rect 302222 212378 302306 212614
rect 302542 212378 302574 212614
rect 301954 212294 302574 212378
rect 301954 212058 301986 212294
rect 302222 212058 302306 212294
rect 302542 212058 302574 212294
rect 301954 176614 302574 212058
rect 301954 176378 301986 176614
rect 302222 176378 302306 176614
rect 302542 176378 302574 176614
rect 301954 176294 302574 176378
rect 301954 176058 301986 176294
rect 302222 176058 302306 176294
rect 302542 176058 302574 176294
rect 301954 140614 302574 176058
rect 301954 140378 301986 140614
rect 302222 140378 302306 140614
rect 302542 140378 302574 140614
rect 301954 140294 302574 140378
rect 301954 140058 301986 140294
rect 302222 140058 302306 140294
rect 302542 140058 302574 140294
rect 301954 104614 302574 140058
rect 301954 104378 301986 104614
rect 302222 104378 302306 104614
rect 302542 104378 302574 104614
rect 301954 104294 302574 104378
rect 301954 104058 301986 104294
rect 302222 104058 302306 104294
rect 302542 104058 302574 104294
rect 301954 68614 302574 104058
rect 301954 68378 301986 68614
rect 302222 68378 302306 68614
rect 302542 68378 302574 68614
rect 301954 68294 302574 68378
rect 301954 68058 301986 68294
rect 302222 68058 302306 68294
rect 302542 68058 302574 68294
rect 301954 32614 302574 68058
rect 301954 32378 301986 32614
rect 302222 32378 302306 32614
rect 302542 32378 302574 32614
rect 301954 32294 302574 32378
rect 301954 32058 301986 32294
rect 302222 32058 302306 32294
rect 302542 32058 302574 32294
rect 298234 -5382 298266 -5146
rect 298502 -5382 298586 -5146
rect 298822 -5382 298854 -5146
rect 298234 -5466 298854 -5382
rect 298234 -5702 298266 -5466
rect 298502 -5702 298586 -5466
rect 298822 -5702 298854 -5466
rect 298234 -5734 298854 -5702
rect 291954 -6342 291986 -6106
rect 292222 -6342 292306 -6106
rect 292542 -6342 292574 -6106
rect 291954 -6426 292574 -6342
rect 291954 -6662 291986 -6426
rect 292222 -6662 292306 -6426
rect 292542 -6662 292574 -6426
rect 291954 -7654 292574 -6662
rect 301954 -7066 302574 32058
rect 304514 706758 305134 707750
rect 304514 706522 304546 706758
rect 304782 706522 304866 706758
rect 305102 706522 305134 706758
rect 304514 706438 305134 706522
rect 304514 706202 304546 706438
rect 304782 706202 304866 706438
rect 305102 706202 305134 706438
rect 304514 691174 305134 706202
rect 304514 690938 304546 691174
rect 304782 690938 304866 691174
rect 305102 690938 305134 691174
rect 304514 690854 305134 690938
rect 304514 690618 304546 690854
rect 304782 690618 304866 690854
rect 305102 690618 305134 690854
rect 304514 655174 305134 690618
rect 304514 654938 304546 655174
rect 304782 654938 304866 655174
rect 305102 654938 305134 655174
rect 304514 654854 305134 654938
rect 304514 654618 304546 654854
rect 304782 654618 304866 654854
rect 305102 654618 305134 654854
rect 304514 619174 305134 654618
rect 304514 618938 304546 619174
rect 304782 618938 304866 619174
rect 305102 618938 305134 619174
rect 304514 618854 305134 618938
rect 304514 618618 304546 618854
rect 304782 618618 304866 618854
rect 305102 618618 305134 618854
rect 304514 583174 305134 618618
rect 304514 582938 304546 583174
rect 304782 582938 304866 583174
rect 305102 582938 305134 583174
rect 304514 582854 305134 582938
rect 304514 582618 304546 582854
rect 304782 582618 304866 582854
rect 305102 582618 305134 582854
rect 304514 547174 305134 582618
rect 304514 546938 304546 547174
rect 304782 546938 304866 547174
rect 305102 546938 305134 547174
rect 304514 546854 305134 546938
rect 304514 546618 304546 546854
rect 304782 546618 304866 546854
rect 305102 546618 305134 546854
rect 304514 511174 305134 546618
rect 304514 510938 304546 511174
rect 304782 510938 304866 511174
rect 305102 510938 305134 511174
rect 304514 510854 305134 510938
rect 304514 510618 304546 510854
rect 304782 510618 304866 510854
rect 305102 510618 305134 510854
rect 304514 475174 305134 510618
rect 304514 474938 304546 475174
rect 304782 474938 304866 475174
rect 305102 474938 305134 475174
rect 304514 474854 305134 474938
rect 304514 474618 304546 474854
rect 304782 474618 304866 474854
rect 305102 474618 305134 474854
rect 304514 439174 305134 474618
rect 304514 438938 304546 439174
rect 304782 438938 304866 439174
rect 305102 438938 305134 439174
rect 304514 438854 305134 438938
rect 304514 438618 304546 438854
rect 304782 438618 304866 438854
rect 305102 438618 305134 438854
rect 304514 403174 305134 438618
rect 304514 402938 304546 403174
rect 304782 402938 304866 403174
rect 305102 402938 305134 403174
rect 304514 402854 305134 402938
rect 304514 402618 304546 402854
rect 304782 402618 304866 402854
rect 305102 402618 305134 402854
rect 304514 367174 305134 402618
rect 304514 366938 304546 367174
rect 304782 366938 304866 367174
rect 305102 366938 305134 367174
rect 304514 366854 305134 366938
rect 304514 366618 304546 366854
rect 304782 366618 304866 366854
rect 305102 366618 305134 366854
rect 304514 331174 305134 366618
rect 304514 330938 304546 331174
rect 304782 330938 304866 331174
rect 305102 330938 305134 331174
rect 304514 330854 305134 330938
rect 304514 330618 304546 330854
rect 304782 330618 304866 330854
rect 305102 330618 305134 330854
rect 304514 295174 305134 330618
rect 304514 294938 304546 295174
rect 304782 294938 304866 295174
rect 305102 294938 305134 295174
rect 304514 294854 305134 294938
rect 304514 294618 304546 294854
rect 304782 294618 304866 294854
rect 305102 294618 305134 294854
rect 304514 259174 305134 294618
rect 304514 258938 304546 259174
rect 304782 258938 304866 259174
rect 305102 258938 305134 259174
rect 304514 258854 305134 258938
rect 304514 258618 304546 258854
rect 304782 258618 304866 258854
rect 305102 258618 305134 258854
rect 304514 223174 305134 258618
rect 304514 222938 304546 223174
rect 304782 222938 304866 223174
rect 305102 222938 305134 223174
rect 304514 222854 305134 222938
rect 304514 222618 304546 222854
rect 304782 222618 304866 222854
rect 305102 222618 305134 222854
rect 304514 187174 305134 222618
rect 304514 186938 304546 187174
rect 304782 186938 304866 187174
rect 305102 186938 305134 187174
rect 304514 186854 305134 186938
rect 304514 186618 304546 186854
rect 304782 186618 304866 186854
rect 305102 186618 305134 186854
rect 304514 151174 305134 186618
rect 304514 150938 304546 151174
rect 304782 150938 304866 151174
rect 305102 150938 305134 151174
rect 304514 150854 305134 150938
rect 304514 150618 304546 150854
rect 304782 150618 304866 150854
rect 305102 150618 305134 150854
rect 304514 115174 305134 150618
rect 304514 114938 304546 115174
rect 304782 114938 304866 115174
rect 305102 114938 305134 115174
rect 304514 114854 305134 114938
rect 304514 114618 304546 114854
rect 304782 114618 304866 114854
rect 305102 114618 305134 114854
rect 304514 79174 305134 114618
rect 304514 78938 304546 79174
rect 304782 78938 304866 79174
rect 305102 78938 305134 79174
rect 304514 78854 305134 78938
rect 304514 78618 304546 78854
rect 304782 78618 304866 78854
rect 305102 78618 305134 78854
rect 304514 43174 305134 78618
rect 304514 42938 304546 43174
rect 304782 42938 304866 43174
rect 305102 42938 305134 43174
rect 304514 42854 305134 42938
rect 304514 42618 304546 42854
rect 304782 42618 304866 42854
rect 305102 42618 305134 42854
rect 304514 7174 305134 42618
rect 304514 6938 304546 7174
rect 304782 6938 304866 7174
rect 305102 6938 305134 7174
rect 304514 6854 305134 6938
rect 304514 6618 304546 6854
rect 304782 6618 304866 6854
rect 305102 6618 305134 6854
rect 304514 -2266 305134 6618
rect 304514 -2502 304546 -2266
rect 304782 -2502 304866 -2266
rect 305102 -2502 305134 -2266
rect 304514 -2586 305134 -2502
rect 304514 -2822 304546 -2586
rect 304782 -2822 304866 -2586
rect 305102 -2822 305134 -2586
rect 304514 -3814 305134 -2822
rect 308234 694894 308854 708122
rect 308234 694658 308266 694894
rect 308502 694658 308586 694894
rect 308822 694658 308854 694894
rect 308234 694574 308854 694658
rect 308234 694338 308266 694574
rect 308502 694338 308586 694574
rect 308822 694338 308854 694574
rect 308234 658894 308854 694338
rect 308234 658658 308266 658894
rect 308502 658658 308586 658894
rect 308822 658658 308854 658894
rect 308234 658574 308854 658658
rect 308234 658338 308266 658574
rect 308502 658338 308586 658574
rect 308822 658338 308854 658574
rect 308234 622894 308854 658338
rect 308234 622658 308266 622894
rect 308502 622658 308586 622894
rect 308822 622658 308854 622894
rect 308234 622574 308854 622658
rect 308234 622338 308266 622574
rect 308502 622338 308586 622574
rect 308822 622338 308854 622574
rect 308234 586894 308854 622338
rect 308234 586658 308266 586894
rect 308502 586658 308586 586894
rect 308822 586658 308854 586894
rect 308234 586574 308854 586658
rect 308234 586338 308266 586574
rect 308502 586338 308586 586574
rect 308822 586338 308854 586574
rect 308234 550894 308854 586338
rect 308234 550658 308266 550894
rect 308502 550658 308586 550894
rect 308822 550658 308854 550894
rect 308234 550574 308854 550658
rect 308234 550338 308266 550574
rect 308502 550338 308586 550574
rect 308822 550338 308854 550574
rect 308234 514894 308854 550338
rect 308234 514658 308266 514894
rect 308502 514658 308586 514894
rect 308822 514658 308854 514894
rect 308234 514574 308854 514658
rect 308234 514338 308266 514574
rect 308502 514338 308586 514574
rect 308822 514338 308854 514574
rect 308234 478894 308854 514338
rect 308234 478658 308266 478894
rect 308502 478658 308586 478894
rect 308822 478658 308854 478894
rect 308234 478574 308854 478658
rect 308234 478338 308266 478574
rect 308502 478338 308586 478574
rect 308822 478338 308854 478574
rect 308234 442894 308854 478338
rect 308234 442658 308266 442894
rect 308502 442658 308586 442894
rect 308822 442658 308854 442894
rect 308234 442574 308854 442658
rect 308234 442338 308266 442574
rect 308502 442338 308586 442574
rect 308822 442338 308854 442574
rect 308234 406894 308854 442338
rect 308234 406658 308266 406894
rect 308502 406658 308586 406894
rect 308822 406658 308854 406894
rect 308234 406574 308854 406658
rect 308234 406338 308266 406574
rect 308502 406338 308586 406574
rect 308822 406338 308854 406574
rect 308234 370894 308854 406338
rect 308234 370658 308266 370894
rect 308502 370658 308586 370894
rect 308822 370658 308854 370894
rect 308234 370574 308854 370658
rect 308234 370338 308266 370574
rect 308502 370338 308586 370574
rect 308822 370338 308854 370574
rect 308234 334894 308854 370338
rect 308234 334658 308266 334894
rect 308502 334658 308586 334894
rect 308822 334658 308854 334894
rect 308234 334574 308854 334658
rect 308234 334338 308266 334574
rect 308502 334338 308586 334574
rect 308822 334338 308854 334574
rect 308234 298894 308854 334338
rect 308234 298658 308266 298894
rect 308502 298658 308586 298894
rect 308822 298658 308854 298894
rect 308234 298574 308854 298658
rect 308234 298338 308266 298574
rect 308502 298338 308586 298574
rect 308822 298338 308854 298574
rect 308234 262894 308854 298338
rect 308234 262658 308266 262894
rect 308502 262658 308586 262894
rect 308822 262658 308854 262894
rect 308234 262574 308854 262658
rect 308234 262338 308266 262574
rect 308502 262338 308586 262574
rect 308822 262338 308854 262574
rect 308234 226894 308854 262338
rect 308234 226658 308266 226894
rect 308502 226658 308586 226894
rect 308822 226658 308854 226894
rect 308234 226574 308854 226658
rect 308234 226338 308266 226574
rect 308502 226338 308586 226574
rect 308822 226338 308854 226574
rect 308234 190894 308854 226338
rect 308234 190658 308266 190894
rect 308502 190658 308586 190894
rect 308822 190658 308854 190894
rect 308234 190574 308854 190658
rect 308234 190338 308266 190574
rect 308502 190338 308586 190574
rect 308822 190338 308854 190574
rect 308234 154894 308854 190338
rect 308234 154658 308266 154894
rect 308502 154658 308586 154894
rect 308822 154658 308854 154894
rect 308234 154574 308854 154658
rect 308234 154338 308266 154574
rect 308502 154338 308586 154574
rect 308822 154338 308854 154574
rect 308234 118894 308854 154338
rect 308234 118658 308266 118894
rect 308502 118658 308586 118894
rect 308822 118658 308854 118894
rect 308234 118574 308854 118658
rect 308234 118338 308266 118574
rect 308502 118338 308586 118574
rect 308822 118338 308854 118574
rect 308234 82894 308854 118338
rect 308234 82658 308266 82894
rect 308502 82658 308586 82894
rect 308822 82658 308854 82894
rect 308234 82574 308854 82658
rect 308234 82338 308266 82574
rect 308502 82338 308586 82574
rect 308822 82338 308854 82574
rect 308234 46894 308854 82338
rect 308234 46658 308266 46894
rect 308502 46658 308586 46894
rect 308822 46658 308854 46894
rect 308234 46574 308854 46658
rect 308234 46338 308266 46574
rect 308502 46338 308586 46574
rect 308822 46338 308854 46574
rect 308234 10894 308854 46338
rect 308234 10658 308266 10894
rect 308502 10658 308586 10894
rect 308822 10658 308854 10894
rect 308234 10574 308854 10658
rect 308234 10338 308266 10574
rect 308502 10338 308586 10574
rect 308822 10338 308854 10574
rect 308234 -4186 308854 10338
rect 310794 705798 311414 705830
rect 310794 705562 310826 705798
rect 311062 705562 311146 705798
rect 311382 705562 311414 705798
rect 310794 705478 311414 705562
rect 310794 705242 310826 705478
rect 311062 705242 311146 705478
rect 311382 705242 311414 705478
rect 310794 669454 311414 705242
rect 310794 669218 310826 669454
rect 311062 669218 311146 669454
rect 311382 669218 311414 669454
rect 310794 669134 311414 669218
rect 310794 668898 310826 669134
rect 311062 668898 311146 669134
rect 311382 668898 311414 669134
rect 310794 633454 311414 668898
rect 310794 633218 310826 633454
rect 311062 633218 311146 633454
rect 311382 633218 311414 633454
rect 310794 633134 311414 633218
rect 310794 632898 310826 633134
rect 311062 632898 311146 633134
rect 311382 632898 311414 633134
rect 310794 597454 311414 632898
rect 310794 597218 310826 597454
rect 311062 597218 311146 597454
rect 311382 597218 311414 597454
rect 310794 597134 311414 597218
rect 310794 596898 310826 597134
rect 311062 596898 311146 597134
rect 311382 596898 311414 597134
rect 310794 561454 311414 596898
rect 310794 561218 310826 561454
rect 311062 561218 311146 561454
rect 311382 561218 311414 561454
rect 310794 561134 311414 561218
rect 310794 560898 310826 561134
rect 311062 560898 311146 561134
rect 311382 560898 311414 561134
rect 310794 525454 311414 560898
rect 310794 525218 310826 525454
rect 311062 525218 311146 525454
rect 311382 525218 311414 525454
rect 310794 525134 311414 525218
rect 310794 524898 310826 525134
rect 311062 524898 311146 525134
rect 311382 524898 311414 525134
rect 310794 489454 311414 524898
rect 310794 489218 310826 489454
rect 311062 489218 311146 489454
rect 311382 489218 311414 489454
rect 310794 489134 311414 489218
rect 310794 488898 310826 489134
rect 311062 488898 311146 489134
rect 311382 488898 311414 489134
rect 310794 453454 311414 488898
rect 310794 453218 310826 453454
rect 311062 453218 311146 453454
rect 311382 453218 311414 453454
rect 310794 453134 311414 453218
rect 310794 452898 310826 453134
rect 311062 452898 311146 453134
rect 311382 452898 311414 453134
rect 310794 417454 311414 452898
rect 310794 417218 310826 417454
rect 311062 417218 311146 417454
rect 311382 417218 311414 417454
rect 310794 417134 311414 417218
rect 310794 416898 310826 417134
rect 311062 416898 311146 417134
rect 311382 416898 311414 417134
rect 310794 381454 311414 416898
rect 310794 381218 310826 381454
rect 311062 381218 311146 381454
rect 311382 381218 311414 381454
rect 310794 381134 311414 381218
rect 310794 380898 310826 381134
rect 311062 380898 311146 381134
rect 311382 380898 311414 381134
rect 310794 345454 311414 380898
rect 310794 345218 310826 345454
rect 311062 345218 311146 345454
rect 311382 345218 311414 345454
rect 310794 345134 311414 345218
rect 310794 344898 310826 345134
rect 311062 344898 311146 345134
rect 311382 344898 311414 345134
rect 310794 309454 311414 344898
rect 310794 309218 310826 309454
rect 311062 309218 311146 309454
rect 311382 309218 311414 309454
rect 310794 309134 311414 309218
rect 310794 308898 310826 309134
rect 311062 308898 311146 309134
rect 311382 308898 311414 309134
rect 310794 273454 311414 308898
rect 310794 273218 310826 273454
rect 311062 273218 311146 273454
rect 311382 273218 311414 273454
rect 310794 273134 311414 273218
rect 310794 272898 310826 273134
rect 311062 272898 311146 273134
rect 311382 272898 311414 273134
rect 310794 237454 311414 272898
rect 310794 237218 310826 237454
rect 311062 237218 311146 237454
rect 311382 237218 311414 237454
rect 310794 237134 311414 237218
rect 310794 236898 310826 237134
rect 311062 236898 311146 237134
rect 311382 236898 311414 237134
rect 310794 201454 311414 236898
rect 310794 201218 310826 201454
rect 311062 201218 311146 201454
rect 311382 201218 311414 201454
rect 310794 201134 311414 201218
rect 310794 200898 310826 201134
rect 311062 200898 311146 201134
rect 311382 200898 311414 201134
rect 310794 165454 311414 200898
rect 310794 165218 310826 165454
rect 311062 165218 311146 165454
rect 311382 165218 311414 165454
rect 310794 165134 311414 165218
rect 310794 164898 310826 165134
rect 311062 164898 311146 165134
rect 311382 164898 311414 165134
rect 310794 129454 311414 164898
rect 310794 129218 310826 129454
rect 311062 129218 311146 129454
rect 311382 129218 311414 129454
rect 310794 129134 311414 129218
rect 310794 128898 310826 129134
rect 311062 128898 311146 129134
rect 311382 128898 311414 129134
rect 310794 93454 311414 128898
rect 310794 93218 310826 93454
rect 311062 93218 311146 93454
rect 311382 93218 311414 93454
rect 310794 93134 311414 93218
rect 310794 92898 310826 93134
rect 311062 92898 311146 93134
rect 311382 92898 311414 93134
rect 310794 57454 311414 92898
rect 310794 57218 310826 57454
rect 311062 57218 311146 57454
rect 311382 57218 311414 57454
rect 310794 57134 311414 57218
rect 310794 56898 310826 57134
rect 311062 56898 311146 57134
rect 311382 56898 311414 57134
rect 310794 21454 311414 56898
rect 310794 21218 310826 21454
rect 311062 21218 311146 21454
rect 311382 21218 311414 21454
rect 310794 21134 311414 21218
rect 310794 20898 310826 21134
rect 311062 20898 311146 21134
rect 311382 20898 311414 21134
rect 310794 -1306 311414 20898
rect 310794 -1542 310826 -1306
rect 311062 -1542 311146 -1306
rect 311382 -1542 311414 -1306
rect 310794 -1626 311414 -1542
rect 310794 -1862 310826 -1626
rect 311062 -1862 311146 -1626
rect 311382 -1862 311414 -1626
rect 310794 -1894 311414 -1862
rect 311954 698614 312574 710042
rect 321954 711558 322574 711590
rect 321954 711322 321986 711558
rect 322222 711322 322306 711558
rect 322542 711322 322574 711558
rect 321954 711238 322574 711322
rect 321954 711002 321986 711238
rect 322222 711002 322306 711238
rect 322542 711002 322574 711238
rect 318234 709638 318854 709670
rect 318234 709402 318266 709638
rect 318502 709402 318586 709638
rect 318822 709402 318854 709638
rect 318234 709318 318854 709402
rect 318234 709082 318266 709318
rect 318502 709082 318586 709318
rect 318822 709082 318854 709318
rect 311954 698378 311986 698614
rect 312222 698378 312306 698614
rect 312542 698378 312574 698614
rect 311954 698294 312574 698378
rect 311954 698058 311986 698294
rect 312222 698058 312306 698294
rect 312542 698058 312574 698294
rect 311954 662614 312574 698058
rect 311954 662378 311986 662614
rect 312222 662378 312306 662614
rect 312542 662378 312574 662614
rect 311954 662294 312574 662378
rect 311954 662058 311986 662294
rect 312222 662058 312306 662294
rect 312542 662058 312574 662294
rect 311954 626614 312574 662058
rect 311954 626378 311986 626614
rect 312222 626378 312306 626614
rect 312542 626378 312574 626614
rect 311954 626294 312574 626378
rect 311954 626058 311986 626294
rect 312222 626058 312306 626294
rect 312542 626058 312574 626294
rect 311954 590614 312574 626058
rect 311954 590378 311986 590614
rect 312222 590378 312306 590614
rect 312542 590378 312574 590614
rect 311954 590294 312574 590378
rect 311954 590058 311986 590294
rect 312222 590058 312306 590294
rect 312542 590058 312574 590294
rect 311954 554614 312574 590058
rect 311954 554378 311986 554614
rect 312222 554378 312306 554614
rect 312542 554378 312574 554614
rect 311954 554294 312574 554378
rect 311954 554058 311986 554294
rect 312222 554058 312306 554294
rect 312542 554058 312574 554294
rect 311954 518614 312574 554058
rect 311954 518378 311986 518614
rect 312222 518378 312306 518614
rect 312542 518378 312574 518614
rect 311954 518294 312574 518378
rect 311954 518058 311986 518294
rect 312222 518058 312306 518294
rect 312542 518058 312574 518294
rect 311954 482614 312574 518058
rect 311954 482378 311986 482614
rect 312222 482378 312306 482614
rect 312542 482378 312574 482614
rect 311954 482294 312574 482378
rect 311954 482058 311986 482294
rect 312222 482058 312306 482294
rect 312542 482058 312574 482294
rect 311954 446614 312574 482058
rect 311954 446378 311986 446614
rect 312222 446378 312306 446614
rect 312542 446378 312574 446614
rect 311954 446294 312574 446378
rect 311954 446058 311986 446294
rect 312222 446058 312306 446294
rect 312542 446058 312574 446294
rect 311954 410614 312574 446058
rect 311954 410378 311986 410614
rect 312222 410378 312306 410614
rect 312542 410378 312574 410614
rect 311954 410294 312574 410378
rect 311954 410058 311986 410294
rect 312222 410058 312306 410294
rect 312542 410058 312574 410294
rect 311954 374614 312574 410058
rect 311954 374378 311986 374614
rect 312222 374378 312306 374614
rect 312542 374378 312574 374614
rect 311954 374294 312574 374378
rect 311954 374058 311986 374294
rect 312222 374058 312306 374294
rect 312542 374058 312574 374294
rect 311954 338614 312574 374058
rect 311954 338378 311986 338614
rect 312222 338378 312306 338614
rect 312542 338378 312574 338614
rect 311954 338294 312574 338378
rect 311954 338058 311986 338294
rect 312222 338058 312306 338294
rect 312542 338058 312574 338294
rect 311954 302614 312574 338058
rect 311954 302378 311986 302614
rect 312222 302378 312306 302614
rect 312542 302378 312574 302614
rect 311954 302294 312574 302378
rect 311954 302058 311986 302294
rect 312222 302058 312306 302294
rect 312542 302058 312574 302294
rect 311954 266614 312574 302058
rect 311954 266378 311986 266614
rect 312222 266378 312306 266614
rect 312542 266378 312574 266614
rect 311954 266294 312574 266378
rect 311954 266058 311986 266294
rect 312222 266058 312306 266294
rect 312542 266058 312574 266294
rect 311954 230614 312574 266058
rect 311954 230378 311986 230614
rect 312222 230378 312306 230614
rect 312542 230378 312574 230614
rect 311954 230294 312574 230378
rect 311954 230058 311986 230294
rect 312222 230058 312306 230294
rect 312542 230058 312574 230294
rect 311954 194614 312574 230058
rect 311954 194378 311986 194614
rect 312222 194378 312306 194614
rect 312542 194378 312574 194614
rect 311954 194294 312574 194378
rect 311954 194058 311986 194294
rect 312222 194058 312306 194294
rect 312542 194058 312574 194294
rect 311954 158614 312574 194058
rect 311954 158378 311986 158614
rect 312222 158378 312306 158614
rect 312542 158378 312574 158614
rect 311954 158294 312574 158378
rect 311954 158058 311986 158294
rect 312222 158058 312306 158294
rect 312542 158058 312574 158294
rect 311954 122614 312574 158058
rect 311954 122378 311986 122614
rect 312222 122378 312306 122614
rect 312542 122378 312574 122614
rect 311954 122294 312574 122378
rect 311954 122058 311986 122294
rect 312222 122058 312306 122294
rect 312542 122058 312574 122294
rect 311954 86614 312574 122058
rect 311954 86378 311986 86614
rect 312222 86378 312306 86614
rect 312542 86378 312574 86614
rect 311954 86294 312574 86378
rect 311954 86058 311986 86294
rect 312222 86058 312306 86294
rect 312542 86058 312574 86294
rect 311954 50614 312574 86058
rect 311954 50378 311986 50614
rect 312222 50378 312306 50614
rect 312542 50378 312574 50614
rect 311954 50294 312574 50378
rect 311954 50058 311986 50294
rect 312222 50058 312306 50294
rect 312542 50058 312574 50294
rect 311954 14614 312574 50058
rect 311954 14378 311986 14614
rect 312222 14378 312306 14614
rect 312542 14378 312574 14614
rect 311954 14294 312574 14378
rect 311954 14058 311986 14294
rect 312222 14058 312306 14294
rect 312542 14058 312574 14294
rect 308234 -4422 308266 -4186
rect 308502 -4422 308586 -4186
rect 308822 -4422 308854 -4186
rect 308234 -4506 308854 -4422
rect 308234 -4742 308266 -4506
rect 308502 -4742 308586 -4506
rect 308822 -4742 308854 -4506
rect 308234 -5734 308854 -4742
rect 301954 -7302 301986 -7066
rect 302222 -7302 302306 -7066
rect 302542 -7302 302574 -7066
rect 301954 -7386 302574 -7302
rect 301954 -7622 301986 -7386
rect 302222 -7622 302306 -7386
rect 302542 -7622 302574 -7386
rect 301954 -7654 302574 -7622
rect 311954 -6106 312574 14058
rect 314514 707718 315134 707750
rect 314514 707482 314546 707718
rect 314782 707482 314866 707718
rect 315102 707482 315134 707718
rect 314514 707398 315134 707482
rect 314514 707162 314546 707398
rect 314782 707162 314866 707398
rect 315102 707162 315134 707398
rect 314514 673174 315134 707162
rect 314514 672938 314546 673174
rect 314782 672938 314866 673174
rect 315102 672938 315134 673174
rect 314514 672854 315134 672938
rect 314514 672618 314546 672854
rect 314782 672618 314866 672854
rect 315102 672618 315134 672854
rect 314514 637174 315134 672618
rect 314514 636938 314546 637174
rect 314782 636938 314866 637174
rect 315102 636938 315134 637174
rect 314514 636854 315134 636938
rect 314514 636618 314546 636854
rect 314782 636618 314866 636854
rect 315102 636618 315134 636854
rect 314514 601174 315134 636618
rect 314514 600938 314546 601174
rect 314782 600938 314866 601174
rect 315102 600938 315134 601174
rect 314514 600854 315134 600938
rect 314514 600618 314546 600854
rect 314782 600618 314866 600854
rect 315102 600618 315134 600854
rect 314514 565174 315134 600618
rect 314514 564938 314546 565174
rect 314782 564938 314866 565174
rect 315102 564938 315134 565174
rect 314514 564854 315134 564938
rect 314514 564618 314546 564854
rect 314782 564618 314866 564854
rect 315102 564618 315134 564854
rect 314514 529174 315134 564618
rect 314514 528938 314546 529174
rect 314782 528938 314866 529174
rect 315102 528938 315134 529174
rect 314514 528854 315134 528938
rect 314514 528618 314546 528854
rect 314782 528618 314866 528854
rect 315102 528618 315134 528854
rect 314514 493174 315134 528618
rect 314514 492938 314546 493174
rect 314782 492938 314866 493174
rect 315102 492938 315134 493174
rect 314514 492854 315134 492938
rect 314514 492618 314546 492854
rect 314782 492618 314866 492854
rect 315102 492618 315134 492854
rect 314514 457174 315134 492618
rect 314514 456938 314546 457174
rect 314782 456938 314866 457174
rect 315102 456938 315134 457174
rect 314514 456854 315134 456938
rect 314514 456618 314546 456854
rect 314782 456618 314866 456854
rect 315102 456618 315134 456854
rect 314514 421174 315134 456618
rect 314514 420938 314546 421174
rect 314782 420938 314866 421174
rect 315102 420938 315134 421174
rect 314514 420854 315134 420938
rect 314514 420618 314546 420854
rect 314782 420618 314866 420854
rect 315102 420618 315134 420854
rect 314514 385174 315134 420618
rect 314514 384938 314546 385174
rect 314782 384938 314866 385174
rect 315102 384938 315134 385174
rect 314514 384854 315134 384938
rect 314514 384618 314546 384854
rect 314782 384618 314866 384854
rect 315102 384618 315134 384854
rect 314514 349174 315134 384618
rect 314514 348938 314546 349174
rect 314782 348938 314866 349174
rect 315102 348938 315134 349174
rect 314514 348854 315134 348938
rect 314514 348618 314546 348854
rect 314782 348618 314866 348854
rect 315102 348618 315134 348854
rect 314514 313174 315134 348618
rect 314514 312938 314546 313174
rect 314782 312938 314866 313174
rect 315102 312938 315134 313174
rect 314514 312854 315134 312938
rect 314514 312618 314546 312854
rect 314782 312618 314866 312854
rect 315102 312618 315134 312854
rect 314514 277174 315134 312618
rect 314514 276938 314546 277174
rect 314782 276938 314866 277174
rect 315102 276938 315134 277174
rect 314514 276854 315134 276938
rect 314514 276618 314546 276854
rect 314782 276618 314866 276854
rect 315102 276618 315134 276854
rect 314514 241174 315134 276618
rect 314514 240938 314546 241174
rect 314782 240938 314866 241174
rect 315102 240938 315134 241174
rect 314514 240854 315134 240938
rect 314514 240618 314546 240854
rect 314782 240618 314866 240854
rect 315102 240618 315134 240854
rect 314514 205174 315134 240618
rect 314514 204938 314546 205174
rect 314782 204938 314866 205174
rect 315102 204938 315134 205174
rect 314514 204854 315134 204938
rect 314514 204618 314546 204854
rect 314782 204618 314866 204854
rect 315102 204618 315134 204854
rect 314514 169174 315134 204618
rect 314514 168938 314546 169174
rect 314782 168938 314866 169174
rect 315102 168938 315134 169174
rect 314514 168854 315134 168938
rect 314514 168618 314546 168854
rect 314782 168618 314866 168854
rect 315102 168618 315134 168854
rect 314514 133174 315134 168618
rect 314514 132938 314546 133174
rect 314782 132938 314866 133174
rect 315102 132938 315134 133174
rect 314514 132854 315134 132938
rect 314514 132618 314546 132854
rect 314782 132618 314866 132854
rect 315102 132618 315134 132854
rect 314514 97174 315134 132618
rect 314514 96938 314546 97174
rect 314782 96938 314866 97174
rect 315102 96938 315134 97174
rect 314514 96854 315134 96938
rect 314514 96618 314546 96854
rect 314782 96618 314866 96854
rect 315102 96618 315134 96854
rect 314514 61174 315134 96618
rect 314514 60938 314546 61174
rect 314782 60938 314866 61174
rect 315102 60938 315134 61174
rect 314514 60854 315134 60938
rect 314514 60618 314546 60854
rect 314782 60618 314866 60854
rect 315102 60618 315134 60854
rect 314514 25174 315134 60618
rect 314514 24938 314546 25174
rect 314782 24938 314866 25174
rect 315102 24938 315134 25174
rect 314514 24854 315134 24938
rect 314514 24618 314546 24854
rect 314782 24618 314866 24854
rect 315102 24618 315134 24854
rect 314514 -3226 315134 24618
rect 314514 -3462 314546 -3226
rect 314782 -3462 314866 -3226
rect 315102 -3462 315134 -3226
rect 314514 -3546 315134 -3462
rect 314514 -3782 314546 -3546
rect 314782 -3782 314866 -3546
rect 315102 -3782 315134 -3546
rect 314514 -3814 315134 -3782
rect 318234 676894 318854 709082
rect 318234 676658 318266 676894
rect 318502 676658 318586 676894
rect 318822 676658 318854 676894
rect 318234 676574 318854 676658
rect 318234 676338 318266 676574
rect 318502 676338 318586 676574
rect 318822 676338 318854 676574
rect 318234 640894 318854 676338
rect 318234 640658 318266 640894
rect 318502 640658 318586 640894
rect 318822 640658 318854 640894
rect 318234 640574 318854 640658
rect 318234 640338 318266 640574
rect 318502 640338 318586 640574
rect 318822 640338 318854 640574
rect 318234 604894 318854 640338
rect 318234 604658 318266 604894
rect 318502 604658 318586 604894
rect 318822 604658 318854 604894
rect 318234 604574 318854 604658
rect 318234 604338 318266 604574
rect 318502 604338 318586 604574
rect 318822 604338 318854 604574
rect 318234 568894 318854 604338
rect 318234 568658 318266 568894
rect 318502 568658 318586 568894
rect 318822 568658 318854 568894
rect 318234 568574 318854 568658
rect 318234 568338 318266 568574
rect 318502 568338 318586 568574
rect 318822 568338 318854 568574
rect 318234 532894 318854 568338
rect 318234 532658 318266 532894
rect 318502 532658 318586 532894
rect 318822 532658 318854 532894
rect 318234 532574 318854 532658
rect 318234 532338 318266 532574
rect 318502 532338 318586 532574
rect 318822 532338 318854 532574
rect 318234 496894 318854 532338
rect 318234 496658 318266 496894
rect 318502 496658 318586 496894
rect 318822 496658 318854 496894
rect 318234 496574 318854 496658
rect 318234 496338 318266 496574
rect 318502 496338 318586 496574
rect 318822 496338 318854 496574
rect 318234 460894 318854 496338
rect 318234 460658 318266 460894
rect 318502 460658 318586 460894
rect 318822 460658 318854 460894
rect 318234 460574 318854 460658
rect 318234 460338 318266 460574
rect 318502 460338 318586 460574
rect 318822 460338 318854 460574
rect 318234 424894 318854 460338
rect 318234 424658 318266 424894
rect 318502 424658 318586 424894
rect 318822 424658 318854 424894
rect 318234 424574 318854 424658
rect 318234 424338 318266 424574
rect 318502 424338 318586 424574
rect 318822 424338 318854 424574
rect 318234 388894 318854 424338
rect 318234 388658 318266 388894
rect 318502 388658 318586 388894
rect 318822 388658 318854 388894
rect 318234 388574 318854 388658
rect 318234 388338 318266 388574
rect 318502 388338 318586 388574
rect 318822 388338 318854 388574
rect 318234 352894 318854 388338
rect 318234 352658 318266 352894
rect 318502 352658 318586 352894
rect 318822 352658 318854 352894
rect 318234 352574 318854 352658
rect 318234 352338 318266 352574
rect 318502 352338 318586 352574
rect 318822 352338 318854 352574
rect 318234 316894 318854 352338
rect 318234 316658 318266 316894
rect 318502 316658 318586 316894
rect 318822 316658 318854 316894
rect 318234 316574 318854 316658
rect 318234 316338 318266 316574
rect 318502 316338 318586 316574
rect 318822 316338 318854 316574
rect 318234 280894 318854 316338
rect 318234 280658 318266 280894
rect 318502 280658 318586 280894
rect 318822 280658 318854 280894
rect 318234 280574 318854 280658
rect 318234 280338 318266 280574
rect 318502 280338 318586 280574
rect 318822 280338 318854 280574
rect 318234 244894 318854 280338
rect 318234 244658 318266 244894
rect 318502 244658 318586 244894
rect 318822 244658 318854 244894
rect 318234 244574 318854 244658
rect 318234 244338 318266 244574
rect 318502 244338 318586 244574
rect 318822 244338 318854 244574
rect 318234 208894 318854 244338
rect 318234 208658 318266 208894
rect 318502 208658 318586 208894
rect 318822 208658 318854 208894
rect 318234 208574 318854 208658
rect 318234 208338 318266 208574
rect 318502 208338 318586 208574
rect 318822 208338 318854 208574
rect 318234 172894 318854 208338
rect 318234 172658 318266 172894
rect 318502 172658 318586 172894
rect 318822 172658 318854 172894
rect 318234 172574 318854 172658
rect 318234 172338 318266 172574
rect 318502 172338 318586 172574
rect 318822 172338 318854 172574
rect 318234 136894 318854 172338
rect 318234 136658 318266 136894
rect 318502 136658 318586 136894
rect 318822 136658 318854 136894
rect 318234 136574 318854 136658
rect 318234 136338 318266 136574
rect 318502 136338 318586 136574
rect 318822 136338 318854 136574
rect 318234 100894 318854 136338
rect 318234 100658 318266 100894
rect 318502 100658 318586 100894
rect 318822 100658 318854 100894
rect 318234 100574 318854 100658
rect 318234 100338 318266 100574
rect 318502 100338 318586 100574
rect 318822 100338 318854 100574
rect 318234 64894 318854 100338
rect 318234 64658 318266 64894
rect 318502 64658 318586 64894
rect 318822 64658 318854 64894
rect 318234 64574 318854 64658
rect 318234 64338 318266 64574
rect 318502 64338 318586 64574
rect 318822 64338 318854 64574
rect 318234 28894 318854 64338
rect 318234 28658 318266 28894
rect 318502 28658 318586 28894
rect 318822 28658 318854 28894
rect 318234 28574 318854 28658
rect 318234 28338 318266 28574
rect 318502 28338 318586 28574
rect 318822 28338 318854 28574
rect 318234 -5146 318854 28338
rect 320794 704838 321414 705830
rect 320794 704602 320826 704838
rect 321062 704602 321146 704838
rect 321382 704602 321414 704838
rect 320794 704518 321414 704602
rect 320794 704282 320826 704518
rect 321062 704282 321146 704518
rect 321382 704282 321414 704518
rect 320794 687454 321414 704282
rect 320794 687218 320826 687454
rect 321062 687218 321146 687454
rect 321382 687218 321414 687454
rect 320794 687134 321414 687218
rect 320794 686898 320826 687134
rect 321062 686898 321146 687134
rect 321382 686898 321414 687134
rect 320794 651454 321414 686898
rect 320794 651218 320826 651454
rect 321062 651218 321146 651454
rect 321382 651218 321414 651454
rect 320794 651134 321414 651218
rect 320794 650898 320826 651134
rect 321062 650898 321146 651134
rect 321382 650898 321414 651134
rect 320794 615454 321414 650898
rect 320794 615218 320826 615454
rect 321062 615218 321146 615454
rect 321382 615218 321414 615454
rect 320794 615134 321414 615218
rect 320794 614898 320826 615134
rect 321062 614898 321146 615134
rect 321382 614898 321414 615134
rect 320794 579454 321414 614898
rect 320794 579218 320826 579454
rect 321062 579218 321146 579454
rect 321382 579218 321414 579454
rect 320794 579134 321414 579218
rect 320794 578898 320826 579134
rect 321062 578898 321146 579134
rect 321382 578898 321414 579134
rect 320794 543454 321414 578898
rect 320794 543218 320826 543454
rect 321062 543218 321146 543454
rect 321382 543218 321414 543454
rect 320794 543134 321414 543218
rect 320794 542898 320826 543134
rect 321062 542898 321146 543134
rect 321382 542898 321414 543134
rect 320794 507454 321414 542898
rect 320794 507218 320826 507454
rect 321062 507218 321146 507454
rect 321382 507218 321414 507454
rect 320794 507134 321414 507218
rect 320794 506898 320826 507134
rect 321062 506898 321146 507134
rect 321382 506898 321414 507134
rect 320794 471454 321414 506898
rect 320794 471218 320826 471454
rect 321062 471218 321146 471454
rect 321382 471218 321414 471454
rect 320794 471134 321414 471218
rect 320794 470898 320826 471134
rect 321062 470898 321146 471134
rect 321382 470898 321414 471134
rect 320794 435454 321414 470898
rect 320794 435218 320826 435454
rect 321062 435218 321146 435454
rect 321382 435218 321414 435454
rect 320794 435134 321414 435218
rect 320794 434898 320826 435134
rect 321062 434898 321146 435134
rect 321382 434898 321414 435134
rect 320794 399454 321414 434898
rect 320794 399218 320826 399454
rect 321062 399218 321146 399454
rect 321382 399218 321414 399454
rect 320794 399134 321414 399218
rect 320794 398898 320826 399134
rect 321062 398898 321146 399134
rect 321382 398898 321414 399134
rect 320794 363454 321414 398898
rect 320794 363218 320826 363454
rect 321062 363218 321146 363454
rect 321382 363218 321414 363454
rect 320794 363134 321414 363218
rect 320794 362898 320826 363134
rect 321062 362898 321146 363134
rect 321382 362898 321414 363134
rect 320794 327454 321414 362898
rect 320794 327218 320826 327454
rect 321062 327218 321146 327454
rect 321382 327218 321414 327454
rect 320794 327134 321414 327218
rect 320794 326898 320826 327134
rect 321062 326898 321146 327134
rect 321382 326898 321414 327134
rect 320794 291454 321414 326898
rect 320794 291218 320826 291454
rect 321062 291218 321146 291454
rect 321382 291218 321414 291454
rect 320794 291134 321414 291218
rect 320794 290898 320826 291134
rect 321062 290898 321146 291134
rect 321382 290898 321414 291134
rect 320794 255454 321414 290898
rect 320794 255218 320826 255454
rect 321062 255218 321146 255454
rect 321382 255218 321414 255454
rect 320794 255134 321414 255218
rect 320794 254898 320826 255134
rect 321062 254898 321146 255134
rect 321382 254898 321414 255134
rect 320794 219454 321414 254898
rect 320794 219218 320826 219454
rect 321062 219218 321146 219454
rect 321382 219218 321414 219454
rect 320794 219134 321414 219218
rect 320794 218898 320826 219134
rect 321062 218898 321146 219134
rect 321382 218898 321414 219134
rect 320794 183454 321414 218898
rect 320794 183218 320826 183454
rect 321062 183218 321146 183454
rect 321382 183218 321414 183454
rect 320794 183134 321414 183218
rect 320794 182898 320826 183134
rect 321062 182898 321146 183134
rect 321382 182898 321414 183134
rect 320794 147454 321414 182898
rect 320794 147218 320826 147454
rect 321062 147218 321146 147454
rect 321382 147218 321414 147454
rect 320794 147134 321414 147218
rect 320794 146898 320826 147134
rect 321062 146898 321146 147134
rect 321382 146898 321414 147134
rect 320794 111454 321414 146898
rect 320794 111218 320826 111454
rect 321062 111218 321146 111454
rect 321382 111218 321414 111454
rect 320794 111134 321414 111218
rect 320794 110898 320826 111134
rect 321062 110898 321146 111134
rect 321382 110898 321414 111134
rect 320794 75454 321414 110898
rect 320794 75218 320826 75454
rect 321062 75218 321146 75454
rect 321382 75218 321414 75454
rect 320794 75134 321414 75218
rect 320794 74898 320826 75134
rect 321062 74898 321146 75134
rect 321382 74898 321414 75134
rect 320794 39454 321414 74898
rect 320794 39218 320826 39454
rect 321062 39218 321146 39454
rect 321382 39218 321414 39454
rect 320794 39134 321414 39218
rect 320794 38898 320826 39134
rect 321062 38898 321146 39134
rect 321382 38898 321414 39134
rect 320794 3454 321414 38898
rect 320794 3218 320826 3454
rect 321062 3218 321146 3454
rect 321382 3218 321414 3454
rect 320794 3134 321414 3218
rect 320794 2898 320826 3134
rect 321062 2898 321146 3134
rect 321382 2898 321414 3134
rect 320794 -346 321414 2898
rect 320794 -582 320826 -346
rect 321062 -582 321146 -346
rect 321382 -582 321414 -346
rect 320794 -666 321414 -582
rect 320794 -902 320826 -666
rect 321062 -902 321146 -666
rect 321382 -902 321414 -666
rect 320794 -1894 321414 -902
rect 321954 680614 322574 711002
rect 331954 710598 332574 711590
rect 331954 710362 331986 710598
rect 332222 710362 332306 710598
rect 332542 710362 332574 710598
rect 331954 710278 332574 710362
rect 331954 710042 331986 710278
rect 332222 710042 332306 710278
rect 332542 710042 332574 710278
rect 328234 708678 328854 709670
rect 328234 708442 328266 708678
rect 328502 708442 328586 708678
rect 328822 708442 328854 708678
rect 328234 708358 328854 708442
rect 328234 708122 328266 708358
rect 328502 708122 328586 708358
rect 328822 708122 328854 708358
rect 321954 680378 321986 680614
rect 322222 680378 322306 680614
rect 322542 680378 322574 680614
rect 321954 680294 322574 680378
rect 321954 680058 321986 680294
rect 322222 680058 322306 680294
rect 322542 680058 322574 680294
rect 321954 644614 322574 680058
rect 321954 644378 321986 644614
rect 322222 644378 322306 644614
rect 322542 644378 322574 644614
rect 321954 644294 322574 644378
rect 321954 644058 321986 644294
rect 322222 644058 322306 644294
rect 322542 644058 322574 644294
rect 321954 608614 322574 644058
rect 321954 608378 321986 608614
rect 322222 608378 322306 608614
rect 322542 608378 322574 608614
rect 321954 608294 322574 608378
rect 321954 608058 321986 608294
rect 322222 608058 322306 608294
rect 322542 608058 322574 608294
rect 321954 572614 322574 608058
rect 321954 572378 321986 572614
rect 322222 572378 322306 572614
rect 322542 572378 322574 572614
rect 321954 572294 322574 572378
rect 321954 572058 321986 572294
rect 322222 572058 322306 572294
rect 322542 572058 322574 572294
rect 321954 536614 322574 572058
rect 321954 536378 321986 536614
rect 322222 536378 322306 536614
rect 322542 536378 322574 536614
rect 321954 536294 322574 536378
rect 321954 536058 321986 536294
rect 322222 536058 322306 536294
rect 322542 536058 322574 536294
rect 321954 500614 322574 536058
rect 321954 500378 321986 500614
rect 322222 500378 322306 500614
rect 322542 500378 322574 500614
rect 321954 500294 322574 500378
rect 321954 500058 321986 500294
rect 322222 500058 322306 500294
rect 322542 500058 322574 500294
rect 321954 464614 322574 500058
rect 321954 464378 321986 464614
rect 322222 464378 322306 464614
rect 322542 464378 322574 464614
rect 321954 464294 322574 464378
rect 321954 464058 321986 464294
rect 322222 464058 322306 464294
rect 322542 464058 322574 464294
rect 321954 428614 322574 464058
rect 321954 428378 321986 428614
rect 322222 428378 322306 428614
rect 322542 428378 322574 428614
rect 321954 428294 322574 428378
rect 321954 428058 321986 428294
rect 322222 428058 322306 428294
rect 322542 428058 322574 428294
rect 321954 392614 322574 428058
rect 321954 392378 321986 392614
rect 322222 392378 322306 392614
rect 322542 392378 322574 392614
rect 321954 392294 322574 392378
rect 321954 392058 321986 392294
rect 322222 392058 322306 392294
rect 322542 392058 322574 392294
rect 321954 356614 322574 392058
rect 321954 356378 321986 356614
rect 322222 356378 322306 356614
rect 322542 356378 322574 356614
rect 321954 356294 322574 356378
rect 321954 356058 321986 356294
rect 322222 356058 322306 356294
rect 322542 356058 322574 356294
rect 321954 320614 322574 356058
rect 321954 320378 321986 320614
rect 322222 320378 322306 320614
rect 322542 320378 322574 320614
rect 321954 320294 322574 320378
rect 321954 320058 321986 320294
rect 322222 320058 322306 320294
rect 322542 320058 322574 320294
rect 321954 284614 322574 320058
rect 321954 284378 321986 284614
rect 322222 284378 322306 284614
rect 322542 284378 322574 284614
rect 321954 284294 322574 284378
rect 321954 284058 321986 284294
rect 322222 284058 322306 284294
rect 322542 284058 322574 284294
rect 321954 248614 322574 284058
rect 321954 248378 321986 248614
rect 322222 248378 322306 248614
rect 322542 248378 322574 248614
rect 321954 248294 322574 248378
rect 321954 248058 321986 248294
rect 322222 248058 322306 248294
rect 322542 248058 322574 248294
rect 321954 212614 322574 248058
rect 321954 212378 321986 212614
rect 322222 212378 322306 212614
rect 322542 212378 322574 212614
rect 321954 212294 322574 212378
rect 321954 212058 321986 212294
rect 322222 212058 322306 212294
rect 322542 212058 322574 212294
rect 321954 176614 322574 212058
rect 321954 176378 321986 176614
rect 322222 176378 322306 176614
rect 322542 176378 322574 176614
rect 321954 176294 322574 176378
rect 321954 176058 321986 176294
rect 322222 176058 322306 176294
rect 322542 176058 322574 176294
rect 321954 140614 322574 176058
rect 321954 140378 321986 140614
rect 322222 140378 322306 140614
rect 322542 140378 322574 140614
rect 321954 140294 322574 140378
rect 321954 140058 321986 140294
rect 322222 140058 322306 140294
rect 322542 140058 322574 140294
rect 321954 104614 322574 140058
rect 321954 104378 321986 104614
rect 322222 104378 322306 104614
rect 322542 104378 322574 104614
rect 321954 104294 322574 104378
rect 321954 104058 321986 104294
rect 322222 104058 322306 104294
rect 322542 104058 322574 104294
rect 321954 68614 322574 104058
rect 321954 68378 321986 68614
rect 322222 68378 322306 68614
rect 322542 68378 322574 68614
rect 321954 68294 322574 68378
rect 321954 68058 321986 68294
rect 322222 68058 322306 68294
rect 322542 68058 322574 68294
rect 321954 32614 322574 68058
rect 321954 32378 321986 32614
rect 322222 32378 322306 32614
rect 322542 32378 322574 32614
rect 321954 32294 322574 32378
rect 321954 32058 321986 32294
rect 322222 32058 322306 32294
rect 322542 32058 322574 32294
rect 318234 -5382 318266 -5146
rect 318502 -5382 318586 -5146
rect 318822 -5382 318854 -5146
rect 318234 -5466 318854 -5382
rect 318234 -5702 318266 -5466
rect 318502 -5702 318586 -5466
rect 318822 -5702 318854 -5466
rect 318234 -5734 318854 -5702
rect 311954 -6342 311986 -6106
rect 312222 -6342 312306 -6106
rect 312542 -6342 312574 -6106
rect 311954 -6426 312574 -6342
rect 311954 -6662 311986 -6426
rect 312222 -6662 312306 -6426
rect 312542 -6662 312574 -6426
rect 311954 -7654 312574 -6662
rect 321954 -7066 322574 32058
rect 324514 706758 325134 707750
rect 324514 706522 324546 706758
rect 324782 706522 324866 706758
rect 325102 706522 325134 706758
rect 324514 706438 325134 706522
rect 324514 706202 324546 706438
rect 324782 706202 324866 706438
rect 325102 706202 325134 706438
rect 324514 691174 325134 706202
rect 324514 690938 324546 691174
rect 324782 690938 324866 691174
rect 325102 690938 325134 691174
rect 324514 690854 325134 690938
rect 324514 690618 324546 690854
rect 324782 690618 324866 690854
rect 325102 690618 325134 690854
rect 324514 655174 325134 690618
rect 324514 654938 324546 655174
rect 324782 654938 324866 655174
rect 325102 654938 325134 655174
rect 324514 654854 325134 654938
rect 324514 654618 324546 654854
rect 324782 654618 324866 654854
rect 325102 654618 325134 654854
rect 324514 619174 325134 654618
rect 324514 618938 324546 619174
rect 324782 618938 324866 619174
rect 325102 618938 325134 619174
rect 324514 618854 325134 618938
rect 324514 618618 324546 618854
rect 324782 618618 324866 618854
rect 325102 618618 325134 618854
rect 324514 583174 325134 618618
rect 324514 582938 324546 583174
rect 324782 582938 324866 583174
rect 325102 582938 325134 583174
rect 324514 582854 325134 582938
rect 324514 582618 324546 582854
rect 324782 582618 324866 582854
rect 325102 582618 325134 582854
rect 324514 547174 325134 582618
rect 324514 546938 324546 547174
rect 324782 546938 324866 547174
rect 325102 546938 325134 547174
rect 324514 546854 325134 546938
rect 324514 546618 324546 546854
rect 324782 546618 324866 546854
rect 325102 546618 325134 546854
rect 324514 511174 325134 546618
rect 324514 510938 324546 511174
rect 324782 510938 324866 511174
rect 325102 510938 325134 511174
rect 324514 510854 325134 510938
rect 324514 510618 324546 510854
rect 324782 510618 324866 510854
rect 325102 510618 325134 510854
rect 324514 475174 325134 510618
rect 324514 474938 324546 475174
rect 324782 474938 324866 475174
rect 325102 474938 325134 475174
rect 324514 474854 325134 474938
rect 324514 474618 324546 474854
rect 324782 474618 324866 474854
rect 325102 474618 325134 474854
rect 324514 439174 325134 474618
rect 324514 438938 324546 439174
rect 324782 438938 324866 439174
rect 325102 438938 325134 439174
rect 324514 438854 325134 438938
rect 324514 438618 324546 438854
rect 324782 438618 324866 438854
rect 325102 438618 325134 438854
rect 324514 403174 325134 438618
rect 324514 402938 324546 403174
rect 324782 402938 324866 403174
rect 325102 402938 325134 403174
rect 324514 402854 325134 402938
rect 324514 402618 324546 402854
rect 324782 402618 324866 402854
rect 325102 402618 325134 402854
rect 324514 367174 325134 402618
rect 324514 366938 324546 367174
rect 324782 366938 324866 367174
rect 325102 366938 325134 367174
rect 324514 366854 325134 366938
rect 324514 366618 324546 366854
rect 324782 366618 324866 366854
rect 325102 366618 325134 366854
rect 324514 331174 325134 366618
rect 324514 330938 324546 331174
rect 324782 330938 324866 331174
rect 325102 330938 325134 331174
rect 324514 330854 325134 330938
rect 324514 330618 324546 330854
rect 324782 330618 324866 330854
rect 325102 330618 325134 330854
rect 324514 295174 325134 330618
rect 324514 294938 324546 295174
rect 324782 294938 324866 295174
rect 325102 294938 325134 295174
rect 324514 294854 325134 294938
rect 324514 294618 324546 294854
rect 324782 294618 324866 294854
rect 325102 294618 325134 294854
rect 324514 259174 325134 294618
rect 324514 258938 324546 259174
rect 324782 258938 324866 259174
rect 325102 258938 325134 259174
rect 324514 258854 325134 258938
rect 324514 258618 324546 258854
rect 324782 258618 324866 258854
rect 325102 258618 325134 258854
rect 324514 223174 325134 258618
rect 324514 222938 324546 223174
rect 324782 222938 324866 223174
rect 325102 222938 325134 223174
rect 324514 222854 325134 222938
rect 324514 222618 324546 222854
rect 324782 222618 324866 222854
rect 325102 222618 325134 222854
rect 324514 187174 325134 222618
rect 324514 186938 324546 187174
rect 324782 186938 324866 187174
rect 325102 186938 325134 187174
rect 324514 186854 325134 186938
rect 324514 186618 324546 186854
rect 324782 186618 324866 186854
rect 325102 186618 325134 186854
rect 324514 151174 325134 186618
rect 324514 150938 324546 151174
rect 324782 150938 324866 151174
rect 325102 150938 325134 151174
rect 324514 150854 325134 150938
rect 324514 150618 324546 150854
rect 324782 150618 324866 150854
rect 325102 150618 325134 150854
rect 324514 115174 325134 150618
rect 324514 114938 324546 115174
rect 324782 114938 324866 115174
rect 325102 114938 325134 115174
rect 324514 114854 325134 114938
rect 324514 114618 324546 114854
rect 324782 114618 324866 114854
rect 325102 114618 325134 114854
rect 324514 79174 325134 114618
rect 324514 78938 324546 79174
rect 324782 78938 324866 79174
rect 325102 78938 325134 79174
rect 324514 78854 325134 78938
rect 324514 78618 324546 78854
rect 324782 78618 324866 78854
rect 325102 78618 325134 78854
rect 324514 43174 325134 78618
rect 324514 42938 324546 43174
rect 324782 42938 324866 43174
rect 325102 42938 325134 43174
rect 324514 42854 325134 42938
rect 324514 42618 324546 42854
rect 324782 42618 324866 42854
rect 325102 42618 325134 42854
rect 324514 7174 325134 42618
rect 324514 6938 324546 7174
rect 324782 6938 324866 7174
rect 325102 6938 325134 7174
rect 324514 6854 325134 6938
rect 324514 6618 324546 6854
rect 324782 6618 324866 6854
rect 325102 6618 325134 6854
rect 324514 -2266 325134 6618
rect 324514 -2502 324546 -2266
rect 324782 -2502 324866 -2266
rect 325102 -2502 325134 -2266
rect 324514 -2586 325134 -2502
rect 324514 -2822 324546 -2586
rect 324782 -2822 324866 -2586
rect 325102 -2822 325134 -2586
rect 324514 -3814 325134 -2822
rect 328234 694894 328854 708122
rect 328234 694658 328266 694894
rect 328502 694658 328586 694894
rect 328822 694658 328854 694894
rect 328234 694574 328854 694658
rect 328234 694338 328266 694574
rect 328502 694338 328586 694574
rect 328822 694338 328854 694574
rect 328234 658894 328854 694338
rect 328234 658658 328266 658894
rect 328502 658658 328586 658894
rect 328822 658658 328854 658894
rect 328234 658574 328854 658658
rect 328234 658338 328266 658574
rect 328502 658338 328586 658574
rect 328822 658338 328854 658574
rect 328234 622894 328854 658338
rect 328234 622658 328266 622894
rect 328502 622658 328586 622894
rect 328822 622658 328854 622894
rect 328234 622574 328854 622658
rect 328234 622338 328266 622574
rect 328502 622338 328586 622574
rect 328822 622338 328854 622574
rect 328234 586894 328854 622338
rect 328234 586658 328266 586894
rect 328502 586658 328586 586894
rect 328822 586658 328854 586894
rect 328234 586574 328854 586658
rect 328234 586338 328266 586574
rect 328502 586338 328586 586574
rect 328822 586338 328854 586574
rect 328234 550894 328854 586338
rect 328234 550658 328266 550894
rect 328502 550658 328586 550894
rect 328822 550658 328854 550894
rect 328234 550574 328854 550658
rect 328234 550338 328266 550574
rect 328502 550338 328586 550574
rect 328822 550338 328854 550574
rect 328234 514894 328854 550338
rect 328234 514658 328266 514894
rect 328502 514658 328586 514894
rect 328822 514658 328854 514894
rect 328234 514574 328854 514658
rect 328234 514338 328266 514574
rect 328502 514338 328586 514574
rect 328822 514338 328854 514574
rect 328234 478894 328854 514338
rect 328234 478658 328266 478894
rect 328502 478658 328586 478894
rect 328822 478658 328854 478894
rect 328234 478574 328854 478658
rect 328234 478338 328266 478574
rect 328502 478338 328586 478574
rect 328822 478338 328854 478574
rect 328234 442894 328854 478338
rect 328234 442658 328266 442894
rect 328502 442658 328586 442894
rect 328822 442658 328854 442894
rect 328234 442574 328854 442658
rect 328234 442338 328266 442574
rect 328502 442338 328586 442574
rect 328822 442338 328854 442574
rect 328234 406894 328854 442338
rect 328234 406658 328266 406894
rect 328502 406658 328586 406894
rect 328822 406658 328854 406894
rect 328234 406574 328854 406658
rect 328234 406338 328266 406574
rect 328502 406338 328586 406574
rect 328822 406338 328854 406574
rect 328234 370894 328854 406338
rect 328234 370658 328266 370894
rect 328502 370658 328586 370894
rect 328822 370658 328854 370894
rect 328234 370574 328854 370658
rect 328234 370338 328266 370574
rect 328502 370338 328586 370574
rect 328822 370338 328854 370574
rect 328234 334894 328854 370338
rect 328234 334658 328266 334894
rect 328502 334658 328586 334894
rect 328822 334658 328854 334894
rect 328234 334574 328854 334658
rect 328234 334338 328266 334574
rect 328502 334338 328586 334574
rect 328822 334338 328854 334574
rect 328234 298894 328854 334338
rect 328234 298658 328266 298894
rect 328502 298658 328586 298894
rect 328822 298658 328854 298894
rect 328234 298574 328854 298658
rect 328234 298338 328266 298574
rect 328502 298338 328586 298574
rect 328822 298338 328854 298574
rect 328234 262894 328854 298338
rect 328234 262658 328266 262894
rect 328502 262658 328586 262894
rect 328822 262658 328854 262894
rect 328234 262574 328854 262658
rect 328234 262338 328266 262574
rect 328502 262338 328586 262574
rect 328822 262338 328854 262574
rect 328234 226894 328854 262338
rect 328234 226658 328266 226894
rect 328502 226658 328586 226894
rect 328822 226658 328854 226894
rect 328234 226574 328854 226658
rect 328234 226338 328266 226574
rect 328502 226338 328586 226574
rect 328822 226338 328854 226574
rect 328234 190894 328854 226338
rect 328234 190658 328266 190894
rect 328502 190658 328586 190894
rect 328822 190658 328854 190894
rect 328234 190574 328854 190658
rect 328234 190338 328266 190574
rect 328502 190338 328586 190574
rect 328822 190338 328854 190574
rect 328234 154894 328854 190338
rect 328234 154658 328266 154894
rect 328502 154658 328586 154894
rect 328822 154658 328854 154894
rect 328234 154574 328854 154658
rect 328234 154338 328266 154574
rect 328502 154338 328586 154574
rect 328822 154338 328854 154574
rect 328234 118894 328854 154338
rect 328234 118658 328266 118894
rect 328502 118658 328586 118894
rect 328822 118658 328854 118894
rect 328234 118574 328854 118658
rect 328234 118338 328266 118574
rect 328502 118338 328586 118574
rect 328822 118338 328854 118574
rect 328234 82894 328854 118338
rect 328234 82658 328266 82894
rect 328502 82658 328586 82894
rect 328822 82658 328854 82894
rect 328234 82574 328854 82658
rect 328234 82338 328266 82574
rect 328502 82338 328586 82574
rect 328822 82338 328854 82574
rect 328234 46894 328854 82338
rect 328234 46658 328266 46894
rect 328502 46658 328586 46894
rect 328822 46658 328854 46894
rect 328234 46574 328854 46658
rect 328234 46338 328266 46574
rect 328502 46338 328586 46574
rect 328822 46338 328854 46574
rect 328234 10894 328854 46338
rect 328234 10658 328266 10894
rect 328502 10658 328586 10894
rect 328822 10658 328854 10894
rect 328234 10574 328854 10658
rect 328234 10338 328266 10574
rect 328502 10338 328586 10574
rect 328822 10338 328854 10574
rect 328234 -4186 328854 10338
rect 330794 705798 331414 705830
rect 330794 705562 330826 705798
rect 331062 705562 331146 705798
rect 331382 705562 331414 705798
rect 330794 705478 331414 705562
rect 330794 705242 330826 705478
rect 331062 705242 331146 705478
rect 331382 705242 331414 705478
rect 330794 669454 331414 705242
rect 330794 669218 330826 669454
rect 331062 669218 331146 669454
rect 331382 669218 331414 669454
rect 330794 669134 331414 669218
rect 330794 668898 330826 669134
rect 331062 668898 331146 669134
rect 331382 668898 331414 669134
rect 330794 633454 331414 668898
rect 330794 633218 330826 633454
rect 331062 633218 331146 633454
rect 331382 633218 331414 633454
rect 330794 633134 331414 633218
rect 330794 632898 330826 633134
rect 331062 632898 331146 633134
rect 331382 632898 331414 633134
rect 330794 597454 331414 632898
rect 330794 597218 330826 597454
rect 331062 597218 331146 597454
rect 331382 597218 331414 597454
rect 330794 597134 331414 597218
rect 330794 596898 330826 597134
rect 331062 596898 331146 597134
rect 331382 596898 331414 597134
rect 330794 561454 331414 596898
rect 330794 561218 330826 561454
rect 331062 561218 331146 561454
rect 331382 561218 331414 561454
rect 330794 561134 331414 561218
rect 330794 560898 330826 561134
rect 331062 560898 331146 561134
rect 331382 560898 331414 561134
rect 330794 525454 331414 560898
rect 330794 525218 330826 525454
rect 331062 525218 331146 525454
rect 331382 525218 331414 525454
rect 330794 525134 331414 525218
rect 330794 524898 330826 525134
rect 331062 524898 331146 525134
rect 331382 524898 331414 525134
rect 330794 489454 331414 524898
rect 330794 489218 330826 489454
rect 331062 489218 331146 489454
rect 331382 489218 331414 489454
rect 330794 489134 331414 489218
rect 330794 488898 330826 489134
rect 331062 488898 331146 489134
rect 331382 488898 331414 489134
rect 330794 453454 331414 488898
rect 330794 453218 330826 453454
rect 331062 453218 331146 453454
rect 331382 453218 331414 453454
rect 330794 453134 331414 453218
rect 330794 452898 330826 453134
rect 331062 452898 331146 453134
rect 331382 452898 331414 453134
rect 330794 417454 331414 452898
rect 330794 417218 330826 417454
rect 331062 417218 331146 417454
rect 331382 417218 331414 417454
rect 330794 417134 331414 417218
rect 330794 416898 330826 417134
rect 331062 416898 331146 417134
rect 331382 416898 331414 417134
rect 330794 381454 331414 416898
rect 330794 381218 330826 381454
rect 331062 381218 331146 381454
rect 331382 381218 331414 381454
rect 330794 381134 331414 381218
rect 330794 380898 330826 381134
rect 331062 380898 331146 381134
rect 331382 380898 331414 381134
rect 330794 345454 331414 380898
rect 330794 345218 330826 345454
rect 331062 345218 331146 345454
rect 331382 345218 331414 345454
rect 330794 345134 331414 345218
rect 330794 344898 330826 345134
rect 331062 344898 331146 345134
rect 331382 344898 331414 345134
rect 330794 309454 331414 344898
rect 330794 309218 330826 309454
rect 331062 309218 331146 309454
rect 331382 309218 331414 309454
rect 330794 309134 331414 309218
rect 330794 308898 330826 309134
rect 331062 308898 331146 309134
rect 331382 308898 331414 309134
rect 330794 273454 331414 308898
rect 330794 273218 330826 273454
rect 331062 273218 331146 273454
rect 331382 273218 331414 273454
rect 330794 273134 331414 273218
rect 330794 272898 330826 273134
rect 331062 272898 331146 273134
rect 331382 272898 331414 273134
rect 330794 237454 331414 272898
rect 330794 237218 330826 237454
rect 331062 237218 331146 237454
rect 331382 237218 331414 237454
rect 330794 237134 331414 237218
rect 330794 236898 330826 237134
rect 331062 236898 331146 237134
rect 331382 236898 331414 237134
rect 330794 201454 331414 236898
rect 330794 201218 330826 201454
rect 331062 201218 331146 201454
rect 331382 201218 331414 201454
rect 330794 201134 331414 201218
rect 330794 200898 330826 201134
rect 331062 200898 331146 201134
rect 331382 200898 331414 201134
rect 330794 165454 331414 200898
rect 330794 165218 330826 165454
rect 331062 165218 331146 165454
rect 331382 165218 331414 165454
rect 330794 165134 331414 165218
rect 330794 164898 330826 165134
rect 331062 164898 331146 165134
rect 331382 164898 331414 165134
rect 330794 129454 331414 164898
rect 330794 129218 330826 129454
rect 331062 129218 331146 129454
rect 331382 129218 331414 129454
rect 330794 129134 331414 129218
rect 330794 128898 330826 129134
rect 331062 128898 331146 129134
rect 331382 128898 331414 129134
rect 330794 93454 331414 128898
rect 330794 93218 330826 93454
rect 331062 93218 331146 93454
rect 331382 93218 331414 93454
rect 330794 93134 331414 93218
rect 330794 92898 330826 93134
rect 331062 92898 331146 93134
rect 331382 92898 331414 93134
rect 330794 57454 331414 92898
rect 330794 57218 330826 57454
rect 331062 57218 331146 57454
rect 331382 57218 331414 57454
rect 330794 57134 331414 57218
rect 330794 56898 330826 57134
rect 331062 56898 331146 57134
rect 331382 56898 331414 57134
rect 330794 21454 331414 56898
rect 330794 21218 330826 21454
rect 331062 21218 331146 21454
rect 331382 21218 331414 21454
rect 330794 21134 331414 21218
rect 330794 20898 330826 21134
rect 331062 20898 331146 21134
rect 331382 20898 331414 21134
rect 330794 -1306 331414 20898
rect 330794 -1542 330826 -1306
rect 331062 -1542 331146 -1306
rect 331382 -1542 331414 -1306
rect 330794 -1626 331414 -1542
rect 330794 -1862 330826 -1626
rect 331062 -1862 331146 -1626
rect 331382 -1862 331414 -1626
rect 330794 -1894 331414 -1862
rect 331954 698614 332574 710042
rect 341954 711558 342574 711590
rect 341954 711322 341986 711558
rect 342222 711322 342306 711558
rect 342542 711322 342574 711558
rect 341954 711238 342574 711322
rect 341954 711002 341986 711238
rect 342222 711002 342306 711238
rect 342542 711002 342574 711238
rect 338234 709638 338854 709670
rect 338234 709402 338266 709638
rect 338502 709402 338586 709638
rect 338822 709402 338854 709638
rect 338234 709318 338854 709402
rect 338234 709082 338266 709318
rect 338502 709082 338586 709318
rect 338822 709082 338854 709318
rect 331954 698378 331986 698614
rect 332222 698378 332306 698614
rect 332542 698378 332574 698614
rect 331954 698294 332574 698378
rect 331954 698058 331986 698294
rect 332222 698058 332306 698294
rect 332542 698058 332574 698294
rect 331954 662614 332574 698058
rect 331954 662378 331986 662614
rect 332222 662378 332306 662614
rect 332542 662378 332574 662614
rect 331954 662294 332574 662378
rect 331954 662058 331986 662294
rect 332222 662058 332306 662294
rect 332542 662058 332574 662294
rect 331954 626614 332574 662058
rect 331954 626378 331986 626614
rect 332222 626378 332306 626614
rect 332542 626378 332574 626614
rect 331954 626294 332574 626378
rect 331954 626058 331986 626294
rect 332222 626058 332306 626294
rect 332542 626058 332574 626294
rect 331954 590614 332574 626058
rect 331954 590378 331986 590614
rect 332222 590378 332306 590614
rect 332542 590378 332574 590614
rect 331954 590294 332574 590378
rect 331954 590058 331986 590294
rect 332222 590058 332306 590294
rect 332542 590058 332574 590294
rect 331954 554614 332574 590058
rect 331954 554378 331986 554614
rect 332222 554378 332306 554614
rect 332542 554378 332574 554614
rect 331954 554294 332574 554378
rect 331954 554058 331986 554294
rect 332222 554058 332306 554294
rect 332542 554058 332574 554294
rect 331954 518614 332574 554058
rect 331954 518378 331986 518614
rect 332222 518378 332306 518614
rect 332542 518378 332574 518614
rect 331954 518294 332574 518378
rect 331954 518058 331986 518294
rect 332222 518058 332306 518294
rect 332542 518058 332574 518294
rect 331954 482614 332574 518058
rect 331954 482378 331986 482614
rect 332222 482378 332306 482614
rect 332542 482378 332574 482614
rect 331954 482294 332574 482378
rect 331954 482058 331986 482294
rect 332222 482058 332306 482294
rect 332542 482058 332574 482294
rect 331954 446614 332574 482058
rect 331954 446378 331986 446614
rect 332222 446378 332306 446614
rect 332542 446378 332574 446614
rect 331954 446294 332574 446378
rect 331954 446058 331986 446294
rect 332222 446058 332306 446294
rect 332542 446058 332574 446294
rect 331954 410614 332574 446058
rect 331954 410378 331986 410614
rect 332222 410378 332306 410614
rect 332542 410378 332574 410614
rect 331954 410294 332574 410378
rect 331954 410058 331986 410294
rect 332222 410058 332306 410294
rect 332542 410058 332574 410294
rect 331954 374614 332574 410058
rect 331954 374378 331986 374614
rect 332222 374378 332306 374614
rect 332542 374378 332574 374614
rect 331954 374294 332574 374378
rect 331954 374058 331986 374294
rect 332222 374058 332306 374294
rect 332542 374058 332574 374294
rect 331954 338614 332574 374058
rect 331954 338378 331986 338614
rect 332222 338378 332306 338614
rect 332542 338378 332574 338614
rect 331954 338294 332574 338378
rect 331954 338058 331986 338294
rect 332222 338058 332306 338294
rect 332542 338058 332574 338294
rect 331954 302614 332574 338058
rect 331954 302378 331986 302614
rect 332222 302378 332306 302614
rect 332542 302378 332574 302614
rect 331954 302294 332574 302378
rect 331954 302058 331986 302294
rect 332222 302058 332306 302294
rect 332542 302058 332574 302294
rect 331954 266614 332574 302058
rect 331954 266378 331986 266614
rect 332222 266378 332306 266614
rect 332542 266378 332574 266614
rect 331954 266294 332574 266378
rect 331954 266058 331986 266294
rect 332222 266058 332306 266294
rect 332542 266058 332574 266294
rect 331954 230614 332574 266058
rect 331954 230378 331986 230614
rect 332222 230378 332306 230614
rect 332542 230378 332574 230614
rect 331954 230294 332574 230378
rect 331954 230058 331986 230294
rect 332222 230058 332306 230294
rect 332542 230058 332574 230294
rect 331954 194614 332574 230058
rect 331954 194378 331986 194614
rect 332222 194378 332306 194614
rect 332542 194378 332574 194614
rect 331954 194294 332574 194378
rect 331954 194058 331986 194294
rect 332222 194058 332306 194294
rect 332542 194058 332574 194294
rect 331954 158614 332574 194058
rect 331954 158378 331986 158614
rect 332222 158378 332306 158614
rect 332542 158378 332574 158614
rect 331954 158294 332574 158378
rect 331954 158058 331986 158294
rect 332222 158058 332306 158294
rect 332542 158058 332574 158294
rect 331954 122614 332574 158058
rect 331954 122378 331986 122614
rect 332222 122378 332306 122614
rect 332542 122378 332574 122614
rect 331954 122294 332574 122378
rect 331954 122058 331986 122294
rect 332222 122058 332306 122294
rect 332542 122058 332574 122294
rect 331954 86614 332574 122058
rect 331954 86378 331986 86614
rect 332222 86378 332306 86614
rect 332542 86378 332574 86614
rect 331954 86294 332574 86378
rect 331954 86058 331986 86294
rect 332222 86058 332306 86294
rect 332542 86058 332574 86294
rect 331954 50614 332574 86058
rect 331954 50378 331986 50614
rect 332222 50378 332306 50614
rect 332542 50378 332574 50614
rect 331954 50294 332574 50378
rect 331954 50058 331986 50294
rect 332222 50058 332306 50294
rect 332542 50058 332574 50294
rect 331954 14614 332574 50058
rect 331954 14378 331986 14614
rect 332222 14378 332306 14614
rect 332542 14378 332574 14614
rect 331954 14294 332574 14378
rect 331954 14058 331986 14294
rect 332222 14058 332306 14294
rect 332542 14058 332574 14294
rect 328234 -4422 328266 -4186
rect 328502 -4422 328586 -4186
rect 328822 -4422 328854 -4186
rect 328234 -4506 328854 -4422
rect 328234 -4742 328266 -4506
rect 328502 -4742 328586 -4506
rect 328822 -4742 328854 -4506
rect 328234 -5734 328854 -4742
rect 321954 -7302 321986 -7066
rect 322222 -7302 322306 -7066
rect 322542 -7302 322574 -7066
rect 321954 -7386 322574 -7302
rect 321954 -7622 321986 -7386
rect 322222 -7622 322306 -7386
rect 322542 -7622 322574 -7386
rect 321954 -7654 322574 -7622
rect 331954 -6106 332574 14058
rect 334514 707718 335134 707750
rect 334514 707482 334546 707718
rect 334782 707482 334866 707718
rect 335102 707482 335134 707718
rect 334514 707398 335134 707482
rect 334514 707162 334546 707398
rect 334782 707162 334866 707398
rect 335102 707162 335134 707398
rect 334514 673174 335134 707162
rect 334514 672938 334546 673174
rect 334782 672938 334866 673174
rect 335102 672938 335134 673174
rect 334514 672854 335134 672938
rect 334514 672618 334546 672854
rect 334782 672618 334866 672854
rect 335102 672618 335134 672854
rect 334514 637174 335134 672618
rect 334514 636938 334546 637174
rect 334782 636938 334866 637174
rect 335102 636938 335134 637174
rect 334514 636854 335134 636938
rect 334514 636618 334546 636854
rect 334782 636618 334866 636854
rect 335102 636618 335134 636854
rect 334514 601174 335134 636618
rect 334514 600938 334546 601174
rect 334782 600938 334866 601174
rect 335102 600938 335134 601174
rect 334514 600854 335134 600938
rect 334514 600618 334546 600854
rect 334782 600618 334866 600854
rect 335102 600618 335134 600854
rect 334514 565174 335134 600618
rect 334514 564938 334546 565174
rect 334782 564938 334866 565174
rect 335102 564938 335134 565174
rect 334514 564854 335134 564938
rect 334514 564618 334546 564854
rect 334782 564618 334866 564854
rect 335102 564618 335134 564854
rect 334514 529174 335134 564618
rect 334514 528938 334546 529174
rect 334782 528938 334866 529174
rect 335102 528938 335134 529174
rect 334514 528854 335134 528938
rect 334514 528618 334546 528854
rect 334782 528618 334866 528854
rect 335102 528618 335134 528854
rect 334514 493174 335134 528618
rect 334514 492938 334546 493174
rect 334782 492938 334866 493174
rect 335102 492938 335134 493174
rect 334514 492854 335134 492938
rect 334514 492618 334546 492854
rect 334782 492618 334866 492854
rect 335102 492618 335134 492854
rect 334514 457174 335134 492618
rect 334514 456938 334546 457174
rect 334782 456938 334866 457174
rect 335102 456938 335134 457174
rect 334514 456854 335134 456938
rect 334514 456618 334546 456854
rect 334782 456618 334866 456854
rect 335102 456618 335134 456854
rect 334514 421174 335134 456618
rect 334514 420938 334546 421174
rect 334782 420938 334866 421174
rect 335102 420938 335134 421174
rect 334514 420854 335134 420938
rect 334514 420618 334546 420854
rect 334782 420618 334866 420854
rect 335102 420618 335134 420854
rect 334514 385174 335134 420618
rect 334514 384938 334546 385174
rect 334782 384938 334866 385174
rect 335102 384938 335134 385174
rect 334514 384854 335134 384938
rect 334514 384618 334546 384854
rect 334782 384618 334866 384854
rect 335102 384618 335134 384854
rect 334514 349174 335134 384618
rect 334514 348938 334546 349174
rect 334782 348938 334866 349174
rect 335102 348938 335134 349174
rect 334514 348854 335134 348938
rect 334514 348618 334546 348854
rect 334782 348618 334866 348854
rect 335102 348618 335134 348854
rect 334514 313174 335134 348618
rect 334514 312938 334546 313174
rect 334782 312938 334866 313174
rect 335102 312938 335134 313174
rect 334514 312854 335134 312938
rect 334514 312618 334546 312854
rect 334782 312618 334866 312854
rect 335102 312618 335134 312854
rect 334514 277174 335134 312618
rect 334514 276938 334546 277174
rect 334782 276938 334866 277174
rect 335102 276938 335134 277174
rect 334514 276854 335134 276938
rect 334514 276618 334546 276854
rect 334782 276618 334866 276854
rect 335102 276618 335134 276854
rect 334514 241174 335134 276618
rect 334514 240938 334546 241174
rect 334782 240938 334866 241174
rect 335102 240938 335134 241174
rect 334514 240854 335134 240938
rect 334514 240618 334546 240854
rect 334782 240618 334866 240854
rect 335102 240618 335134 240854
rect 334514 205174 335134 240618
rect 334514 204938 334546 205174
rect 334782 204938 334866 205174
rect 335102 204938 335134 205174
rect 334514 204854 335134 204938
rect 334514 204618 334546 204854
rect 334782 204618 334866 204854
rect 335102 204618 335134 204854
rect 334514 169174 335134 204618
rect 334514 168938 334546 169174
rect 334782 168938 334866 169174
rect 335102 168938 335134 169174
rect 334514 168854 335134 168938
rect 334514 168618 334546 168854
rect 334782 168618 334866 168854
rect 335102 168618 335134 168854
rect 334514 133174 335134 168618
rect 334514 132938 334546 133174
rect 334782 132938 334866 133174
rect 335102 132938 335134 133174
rect 334514 132854 335134 132938
rect 334514 132618 334546 132854
rect 334782 132618 334866 132854
rect 335102 132618 335134 132854
rect 334514 97174 335134 132618
rect 334514 96938 334546 97174
rect 334782 96938 334866 97174
rect 335102 96938 335134 97174
rect 334514 96854 335134 96938
rect 334514 96618 334546 96854
rect 334782 96618 334866 96854
rect 335102 96618 335134 96854
rect 334514 61174 335134 96618
rect 334514 60938 334546 61174
rect 334782 60938 334866 61174
rect 335102 60938 335134 61174
rect 334514 60854 335134 60938
rect 334514 60618 334546 60854
rect 334782 60618 334866 60854
rect 335102 60618 335134 60854
rect 334514 25174 335134 60618
rect 334514 24938 334546 25174
rect 334782 24938 334866 25174
rect 335102 24938 335134 25174
rect 334514 24854 335134 24938
rect 334514 24618 334546 24854
rect 334782 24618 334866 24854
rect 335102 24618 335134 24854
rect 334514 -3226 335134 24618
rect 334514 -3462 334546 -3226
rect 334782 -3462 334866 -3226
rect 335102 -3462 335134 -3226
rect 334514 -3546 335134 -3462
rect 334514 -3782 334546 -3546
rect 334782 -3782 334866 -3546
rect 335102 -3782 335134 -3546
rect 334514 -3814 335134 -3782
rect 338234 676894 338854 709082
rect 338234 676658 338266 676894
rect 338502 676658 338586 676894
rect 338822 676658 338854 676894
rect 338234 676574 338854 676658
rect 338234 676338 338266 676574
rect 338502 676338 338586 676574
rect 338822 676338 338854 676574
rect 338234 640894 338854 676338
rect 338234 640658 338266 640894
rect 338502 640658 338586 640894
rect 338822 640658 338854 640894
rect 338234 640574 338854 640658
rect 338234 640338 338266 640574
rect 338502 640338 338586 640574
rect 338822 640338 338854 640574
rect 338234 604894 338854 640338
rect 338234 604658 338266 604894
rect 338502 604658 338586 604894
rect 338822 604658 338854 604894
rect 338234 604574 338854 604658
rect 338234 604338 338266 604574
rect 338502 604338 338586 604574
rect 338822 604338 338854 604574
rect 338234 568894 338854 604338
rect 338234 568658 338266 568894
rect 338502 568658 338586 568894
rect 338822 568658 338854 568894
rect 338234 568574 338854 568658
rect 338234 568338 338266 568574
rect 338502 568338 338586 568574
rect 338822 568338 338854 568574
rect 338234 532894 338854 568338
rect 338234 532658 338266 532894
rect 338502 532658 338586 532894
rect 338822 532658 338854 532894
rect 338234 532574 338854 532658
rect 338234 532338 338266 532574
rect 338502 532338 338586 532574
rect 338822 532338 338854 532574
rect 338234 496894 338854 532338
rect 338234 496658 338266 496894
rect 338502 496658 338586 496894
rect 338822 496658 338854 496894
rect 338234 496574 338854 496658
rect 338234 496338 338266 496574
rect 338502 496338 338586 496574
rect 338822 496338 338854 496574
rect 338234 460894 338854 496338
rect 338234 460658 338266 460894
rect 338502 460658 338586 460894
rect 338822 460658 338854 460894
rect 338234 460574 338854 460658
rect 338234 460338 338266 460574
rect 338502 460338 338586 460574
rect 338822 460338 338854 460574
rect 338234 424894 338854 460338
rect 338234 424658 338266 424894
rect 338502 424658 338586 424894
rect 338822 424658 338854 424894
rect 338234 424574 338854 424658
rect 338234 424338 338266 424574
rect 338502 424338 338586 424574
rect 338822 424338 338854 424574
rect 338234 388894 338854 424338
rect 338234 388658 338266 388894
rect 338502 388658 338586 388894
rect 338822 388658 338854 388894
rect 338234 388574 338854 388658
rect 338234 388338 338266 388574
rect 338502 388338 338586 388574
rect 338822 388338 338854 388574
rect 338234 352894 338854 388338
rect 338234 352658 338266 352894
rect 338502 352658 338586 352894
rect 338822 352658 338854 352894
rect 338234 352574 338854 352658
rect 338234 352338 338266 352574
rect 338502 352338 338586 352574
rect 338822 352338 338854 352574
rect 338234 316894 338854 352338
rect 338234 316658 338266 316894
rect 338502 316658 338586 316894
rect 338822 316658 338854 316894
rect 338234 316574 338854 316658
rect 338234 316338 338266 316574
rect 338502 316338 338586 316574
rect 338822 316338 338854 316574
rect 338234 280894 338854 316338
rect 338234 280658 338266 280894
rect 338502 280658 338586 280894
rect 338822 280658 338854 280894
rect 338234 280574 338854 280658
rect 338234 280338 338266 280574
rect 338502 280338 338586 280574
rect 338822 280338 338854 280574
rect 338234 244894 338854 280338
rect 338234 244658 338266 244894
rect 338502 244658 338586 244894
rect 338822 244658 338854 244894
rect 338234 244574 338854 244658
rect 338234 244338 338266 244574
rect 338502 244338 338586 244574
rect 338822 244338 338854 244574
rect 338234 208894 338854 244338
rect 338234 208658 338266 208894
rect 338502 208658 338586 208894
rect 338822 208658 338854 208894
rect 338234 208574 338854 208658
rect 338234 208338 338266 208574
rect 338502 208338 338586 208574
rect 338822 208338 338854 208574
rect 338234 172894 338854 208338
rect 338234 172658 338266 172894
rect 338502 172658 338586 172894
rect 338822 172658 338854 172894
rect 338234 172574 338854 172658
rect 338234 172338 338266 172574
rect 338502 172338 338586 172574
rect 338822 172338 338854 172574
rect 338234 136894 338854 172338
rect 338234 136658 338266 136894
rect 338502 136658 338586 136894
rect 338822 136658 338854 136894
rect 338234 136574 338854 136658
rect 338234 136338 338266 136574
rect 338502 136338 338586 136574
rect 338822 136338 338854 136574
rect 338234 100894 338854 136338
rect 338234 100658 338266 100894
rect 338502 100658 338586 100894
rect 338822 100658 338854 100894
rect 338234 100574 338854 100658
rect 338234 100338 338266 100574
rect 338502 100338 338586 100574
rect 338822 100338 338854 100574
rect 338234 64894 338854 100338
rect 338234 64658 338266 64894
rect 338502 64658 338586 64894
rect 338822 64658 338854 64894
rect 338234 64574 338854 64658
rect 338234 64338 338266 64574
rect 338502 64338 338586 64574
rect 338822 64338 338854 64574
rect 338234 28894 338854 64338
rect 338234 28658 338266 28894
rect 338502 28658 338586 28894
rect 338822 28658 338854 28894
rect 338234 28574 338854 28658
rect 338234 28338 338266 28574
rect 338502 28338 338586 28574
rect 338822 28338 338854 28574
rect 338234 -5146 338854 28338
rect 340794 704838 341414 705830
rect 340794 704602 340826 704838
rect 341062 704602 341146 704838
rect 341382 704602 341414 704838
rect 340794 704518 341414 704602
rect 340794 704282 340826 704518
rect 341062 704282 341146 704518
rect 341382 704282 341414 704518
rect 340794 687454 341414 704282
rect 340794 687218 340826 687454
rect 341062 687218 341146 687454
rect 341382 687218 341414 687454
rect 340794 687134 341414 687218
rect 340794 686898 340826 687134
rect 341062 686898 341146 687134
rect 341382 686898 341414 687134
rect 340794 651454 341414 686898
rect 340794 651218 340826 651454
rect 341062 651218 341146 651454
rect 341382 651218 341414 651454
rect 340794 651134 341414 651218
rect 340794 650898 340826 651134
rect 341062 650898 341146 651134
rect 341382 650898 341414 651134
rect 340794 615454 341414 650898
rect 340794 615218 340826 615454
rect 341062 615218 341146 615454
rect 341382 615218 341414 615454
rect 340794 615134 341414 615218
rect 340794 614898 340826 615134
rect 341062 614898 341146 615134
rect 341382 614898 341414 615134
rect 340794 579454 341414 614898
rect 340794 579218 340826 579454
rect 341062 579218 341146 579454
rect 341382 579218 341414 579454
rect 340794 579134 341414 579218
rect 340794 578898 340826 579134
rect 341062 578898 341146 579134
rect 341382 578898 341414 579134
rect 340794 543454 341414 578898
rect 340794 543218 340826 543454
rect 341062 543218 341146 543454
rect 341382 543218 341414 543454
rect 340794 543134 341414 543218
rect 340794 542898 340826 543134
rect 341062 542898 341146 543134
rect 341382 542898 341414 543134
rect 340794 507454 341414 542898
rect 340794 507218 340826 507454
rect 341062 507218 341146 507454
rect 341382 507218 341414 507454
rect 340794 507134 341414 507218
rect 340794 506898 340826 507134
rect 341062 506898 341146 507134
rect 341382 506898 341414 507134
rect 340794 471454 341414 506898
rect 340794 471218 340826 471454
rect 341062 471218 341146 471454
rect 341382 471218 341414 471454
rect 340794 471134 341414 471218
rect 340794 470898 340826 471134
rect 341062 470898 341146 471134
rect 341382 470898 341414 471134
rect 340794 435454 341414 470898
rect 340794 435218 340826 435454
rect 341062 435218 341146 435454
rect 341382 435218 341414 435454
rect 340794 435134 341414 435218
rect 340794 434898 340826 435134
rect 341062 434898 341146 435134
rect 341382 434898 341414 435134
rect 340794 399454 341414 434898
rect 340794 399218 340826 399454
rect 341062 399218 341146 399454
rect 341382 399218 341414 399454
rect 340794 399134 341414 399218
rect 340794 398898 340826 399134
rect 341062 398898 341146 399134
rect 341382 398898 341414 399134
rect 340794 363454 341414 398898
rect 340794 363218 340826 363454
rect 341062 363218 341146 363454
rect 341382 363218 341414 363454
rect 340794 363134 341414 363218
rect 340794 362898 340826 363134
rect 341062 362898 341146 363134
rect 341382 362898 341414 363134
rect 340794 327454 341414 362898
rect 340794 327218 340826 327454
rect 341062 327218 341146 327454
rect 341382 327218 341414 327454
rect 340794 327134 341414 327218
rect 340794 326898 340826 327134
rect 341062 326898 341146 327134
rect 341382 326898 341414 327134
rect 340794 291454 341414 326898
rect 340794 291218 340826 291454
rect 341062 291218 341146 291454
rect 341382 291218 341414 291454
rect 340794 291134 341414 291218
rect 340794 290898 340826 291134
rect 341062 290898 341146 291134
rect 341382 290898 341414 291134
rect 340794 255454 341414 290898
rect 340794 255218 340826 255454
rect 341062 255218 341146 255454
rect 341382 255218 341414 255454
rect 340794 255134 341414 255218
rect 340794 254898 340826 255134
rect 341062 254898 341146 255134
rect 341382 254898 341414 255134
rect 340794 219454 341414 254898
rect 340794 219218 340826 219454
rect 341062 219218 341146 219454
rect 341382 219218 341414 219454
rect 340794 219134 341414 219218
rect 340794 218898 340826 219134
rect 341062 218898 341146 219134
rect 341382 218898 341414 219134
rect 340794 183454 341414 218898
rect 340794 183218 340826 183454
rect 341062 183218 341146 183454
rect 341382 183218 341414 183454
rect 340794 183134 341414 183218
rect 340794 182898 340826 183134
rect 341062 182898 341146 183134
rect 341382 182898 341414 183134
rect 340794 147454 341414 182898
rect 340794 147218 340826 147454
rect 341062 147218 341146 147454
rect 341382 147218 341414 147454
rect 340794 147134 341414 147218
rect 340794 146898 340826 147134
rect 341062 146898 341146 147134
rect 341382 146898 341414 147134
rect 340794 111454 341414 146898
rect 340794 111218 340826 111454
rect 341062 111218 341146 111454
rect 341382 111218 341414 111454
rect 340794 111134 341414 111218
rect 340794 110898 340826 111134
rect 341062 110898 341146 111134
rect 341382 110898 341414 111134
rect 340794 75454 341414 110898
rect 340794 75218 340826 75454
rect 341062 75218 341146 75454
rect 341382 75218 341414 75454
rect 340794 75134 341414 75218
rect 340794 74898 340826 75134
rect 341062 74898 341146 75134
rect 341382 74898 341414 75134
rect 340794 39454 341414 74898
rect 340794 39218 340826 39454
rect 341062 39218 341146 39454
rect 341382 39218 341414 39454
rect 340794 39134 341414 39218
rect 340794 38898 340826 39134
rect 341062 38898 341146 39134
rect 341382 38898 341414 39134
rect 340794 3454 341414 38898
rect 340794 3218 340826 3454
rect 341062 3218 341146 3454
rect 341382 3218 341414 3454
rect 340794 3134 341414 3218
rect 340794 2898 340826 3134
rect 341062 2898 341146 3134
rect 341382 2898 341414 3134
rect 340794 -346 341414 2898
rect 340794 -582 340826 -346
rect 341062 -582 341146 -346
rect 341382 -582 341414 -346
rect 340794 -666 341414 -582
rect 340794 -902 340826 -666
rect 341062 -902 341146 -666
rect 341382 -902 341414 -666
rect 340794 -1894 341414 -902
rect 341954 680614 342574 711002
rect 351954 710598 352574 711590
rect 351954 710362 351986 710598
rect 352222 710362 352306 710598
rect 352542 710362 352574 710598
rect 351954 710278 352574 710362
rect 351954 710042 351986 710278
rect 352222 710042 352306 710278
rect 352542 710042 352574 710278
rect 348234 708678 348854 709670
rect 348234 708442 348266 708678
rect 348502 708442 348586 708678
rect 348822 708442 348854 708678
rect 348234 708358 348854 708442
rect 348234 708122 348266 708358
rect 348502 708122 348586 708358
rect 348822 708122 348854 708358
rect 341954 680378 341986 680614
rect 342222 680378 342306 680614
rect 342542 680378 342574 680614
rect 341954 680294 342574 680378
rect 341954 680058 341986 680294
rect 342222 680058 342306 680294
rect 342542 680058 342574 680294
rect 341954 644614 342574 680058
rect 341954 644378 341986 644614
rect 342222 644378 342306 644614
rect 342542 644378 342574 644614
rect 341954 644294 342574 644378
rect 341954 644058 341986 644294
rect 342222 644058 342306 644294
rect 342542 644058 342574 644294
rect 341954 608614 342574 644058
rect 341954 608378 341986 608614
rect 342222 608378 342306 608614
rect 342542 608378 342574 608614
rect 341954 608294 342574 608378
rect 341954 608058 341986 608294
rect 342222 608058 342306 608294
rect 342542 608058 342574 608294
rect 341954 572614 342574 608058
rect 341954 572378 341986 572614
rect 342222 572378 342306 572614
rect 342542 572378 342574 572614
rect 341954 572294 342574 572378
rect 341954 572058 341986 572294
rect 342222 572058 342306 572294
rect 342542 572058 342574 572294
rect 341954 536614 342574 572058
rect 341954 536378 341986 536614
rect 342222 536378 342306 536614
rect 342542 536378 342574 536614
rect 341954 536294 342574 536378
rect 341954 536058 341986 536294
rect 342222 536058 342306 536294
rect 342542 536058 342574 536294
rect 341954 500614 342574 536058
rect 341954 500378 341986 500614
rect 342222 500378 342306 500614
rect 342542 500378 342574 500614
rect 341954 500294 342574 500378
rect 341954 500058 341986 500294
rect 342222 500058 342306 500294
rect 342542 500058 342574 500294
rect 341954 464614 342574 500058
rect 341954 464378 341986 464614
rect 342222 464378 342306 464614
rect 342542 464378 342574 464614
rect 341954 464294 342574 464378
rect 341954 464058 341986 464294
rect 342222 464058 342306 464294
rect 342542 464058 342574 464294
rect 341954 428614 342574 464058
rect 341954 428378 341986 428614
rect 342222 428378 342306 428614
rect 342542 428378 342574 428614
rect 341954 428294 342574 428378
rect 341954 428058 341986 428294
rect 342222 428058 342306 428294
rect 342542 428058 342574 428294
rect 341954 392614 342574 428058
rect 341954 392378 341986 392614
rect 342222 392378 342306 392614
rect 342542 392378 342574 392614
rect 341954 392294 342574 392378
rect 341954 392058 341986 392294
rect 342222 392058 342306 392294
rect 342542 392058 342574 392294
rect 341954 356614 342574 392058
rect 341954 356378 341986 356614
rect 342222 356378 342306 356614
rect 342542 356378 342574 356614
rect 341954 356294 342574 356378
rect 341954 356058 341986 356294
rect 342222 356058 342306 356294
rect 342542 356058 342574 356294
rect 341954 320614 342574 356058
rect 341954 320378 341986 320614
rect 342222 320378 342306 320614
rect 342542 320378 342574 320614
rect 341954 320294 342574 320378
rect 341954 320058 341986 320294
rect 342222 320058 342306 320294
rect 342542 320058 342574 320294
rect 341954 284614 342574 320058
rect 341954 284378 341986 284614
rect 342222 284378 342306 284614
rect 342542 284378 342574 284614
rect 341954 284294 342574 284378
rect 341954 284058 341986 284294
rect 342222 284058 342306 284294
rect 342542 284058 342574 284294
rect 341954 248614 342574 284058
rect 341954 248378 341986 248614
rect 342222 248378 342306 248614
rect 342542 248378 342574 248614
rect 341954 248294 342574 248378
rect 341954 248058 341986 248294
rect 342222 248058 342306 248294
rect 342542 248058 342574 248294
rect 341954 212614 342574 248058
rect 341954 212378 341986 212614
rect 342222 212378 342306 212614
rect 342542 212378 342574 212614
rect 341954 212294 342574 212378
rect 341954 212058 341986 212294
rect 342222 212058 342306 212294
rect 342542 212058 342574 212294
rect 341954 176614 342574 212058
rect 341954 176378 341986 176614
rect 342222 176378 342306 176614
rect 342542 176378 342574 176614
rect 341954 176294 342574 176378
rect 341954 176058 341986 176294
rect 342222 176058 342306 176294
rect 342542 176058 342574 176294
rect 341954 140614 342574 176058
rect 341954 140378 341986 140614
rect 342222 140378 342306 140614
rect 342542 140378 342574 140614
rect 341954 140294 342574 140378
rect 341954 140058 341986 140294
rect 342222 140058 342306 140294
rect 342542 140058 342574 140294
rect 341954 104614 342574 140058
rect 341954 104378 341986 104614
rect 342222 104378 342306 104614
rect 342542 104378 342574 104614
rect 341954 104294 342574 104378
rect 341954 104058 341986 104294
rect 342222 104058 342306 104294
rect 342542 104058 342574 104294
rect 341954 68614 342574 104058
rect 341954 68378 341986 68614
rect 342222 68378 342306 68614
rect 342542 68378 342574 68614
rect 341954 68294 342574 68378
rect 341954 68058 341986 68294
rect 342222 68058 342306 68294
rect 342542 68058 342574 68294
rect 341954 32614 342574 68058
rect 341954 32378 341986 32614
rect 342222 32378 342306 32614
rect 342542 32378 342574 32614
rect 341954 32294 342574 32378
rect 341954 32058 341986 32294
rect 342222 32058 342306 32294
rect 342542 32058 342574 32294
rect 338234 -5382 338266 -5146
rect 338502 -5382 338586 -5146
rect 338822 -5382 338854 -5146
rect 338234 -5466 338854 -5382
rect 338234 -5702 338266 -5466
rect 338502 -5702 338586 -5466
rect 338822 -5702 338854 -5466
rect 338234 -5734 338854 -5702
rect 331954 -6342 331986 -6106
rect 332222 -6342 332306 -6106
rect 332542 -6342 332574 -6106
rect 331954 -6426 332574 -6342
rect 331954 -6662 331986 -6426
rect 332222 -6662 332306 -6426
rect 332542 -6662 332574 -6426
rect 331954 -7654 332574 -6662
rect 341954 -7066 342574 32058
rect 344514 706758 345134 707750
rect 344514 706522 344546 706758
rect 344782 706522 344866 706758
rect 345102 706522 345134 706758
rect 344514 706438 345134 706522
rect 344514 706202 344546 706438
rect 344782 706202 344866 706438
rect 345102 706202 345134 706438
rect 344514 691174 345134 706202
rect 344514 690938 344546 691174
rect 344782 690938 344866 691174
rect 345102 690938 345134 691174
rect 344514 690854 345134 690938
rect 344514 690618 344546 690854
rect 344782 690618 344866 690854
rect 345102 690618 345134 690854
rect 344514 655174 345134 690618
rect 344514 654938 344546 655174
rect 344782 654938 344866 655174
rect 345102 654938 345134 655174
rect 344514 654854 345134 654938
rect 344514 654618 344546 654854
rect 344782 654618 344866 654854
rect 345102 654618 345134 654854
rect 344514 619174 345134 654618
rect 344514 618938 344546 619174
rect 344782 618938 344866 619174
rect 345102 618938 345134 619174
rect 344514 618854 345134 618938
rect 344514 618618 344546 618854
rect 344782 618618 344866 618854
rect 345102 618618 345134 618854
rect 344514 583174 345134 618618
rect 344514 582938 344546 583174
rect 344782 582938 344866 583174
rect 345102 582938 345134 583174
rect 344514 582854 345134 582938
rect 344514 582618 344546 582854
rect 344782 582618 344866 582854
rect 345102 582618 345134 582854
rect 344514 547174 345134 582618
rect 344514 546938 344546 547174
rect 344782 546938 344866 547174
rect 345102 546938 345134 547174
rect 344514 546854 345134 546938
rect 344514 546618 344546 546854
rect 344782 546618 344866 546854
rect 345102 546618 345134 546854
rect 344514 511174 345134 546618
rect 344514 510938 344546 511174
rect 344782 510938 344866 511174
rect 345102 510938 345134 511174
rect 344514 510854 345134 510938
rect 344514 510618 344546 510854
rect 344782 510618 344866 510854
rect 345102 510618 345134 510854
rect 344514 475174 345134 510618
rect 344514 474938 344546 475174
rect 344782 474938 344866 475174
rect 345102 474938 345134 475174
rect 344514 474854 345134 474938
rect 344514 474618 344546 474854
rect 344782 474618 344866 474854
rect 345102 474618 345134 474854
rect 344514 439174 345134 474618
rect 344514 438938 344546 439174
rect 344782 438938 344866 439174
rect 345102 438938 345134 439174
rect 344514 438854 345134 438938
rect 344514 438618 344546 438854
rect 344782 438618 344866 438854
rect 345102 438618 345134 438854
rect 344514 403174 345134 438618
rect 344514 402938 344546 403174
rect 344782 402938 344866 403174
rect 345102 402938 345134 403174
rect 344514 402854 345134 402938
rect 344514 402618 344546 402854
rect 344782 402618 344866 402854
rect 345102 402618 345134 402854
rect 344514 367174 345134 402618
rect 344514 366938 344546 367174
rect 344782 366938 344866 367174
rect 345102 366938 345134 367174
rect 344514 366854 345134 366938
rect 344514 366618 344546 366854
rect 344782 366618 344866 366854
rect 345102 366618 345134 366854
rect 344514 331174 345134 366618
rect 344514 330938 344546 331174
rect 344782 330938 344866 331174
rect 345102 330938 345134 331174
rect 344514 330854 345134 330938
rect 344514 330618 344546 330854
rect 344782 330618 344866 330854
rect 345102 330618 345134 330854
rect 344514 295174 345134 330618
rect 344514 294938 344546 295174
rect 344782 294938 344866 295174
rect 345102 294938 345134 295174
rect 344514 294854 345134 294938
rect 344514 294618 344546 294854
rect 344782 294618 344866 294854
rect 345102 294618 345134 294854
rect 344514 259174 345134 294618
rect 344514 258938 344546 259174
rect 344782 258938 344866 259174
rect 345102 258938 345134 259174
rect 344514 258854 345134 258938
rect 344514 258618 344546 258854
rect 344782 258618 344866 258854
rect 345102 258618 345134 258854
rect 344514 223174 345134 258618
rect 344514 222938 344546 223174
rect 344782 222938 344866 223174
rect 345102 222938 345134 223174
rect 344514 222854 345134 222938
rect 344514 222618 344546 222854
rect 344782 222618 344866 222854
rect 345102 222618 345134 222854
rect 344514 187174 345134 222618
rect 344514 186938 344546 187174
rect 344782 186938 344866 187174
rect 345102 186938 345134 187174
rect 344514 186854 345134 186938
rect 344514 186618 344546 186854
rect 344782 186618 344866 186854
rect 345102 186618 345134 186854
rect 344514 151174 345134 186618
rect 344514 150938 344546 151174
rect 344782 150938 344866 151174
rect 345102 150938 345134 151174
rect 344514 150854 345134 150938
rect 344514 150618 344546 150854
rect 344782 150618 344866 150854
rect 345102 150618 345134 150854
rect 344514 115174 345134 150618
rect 344514 114938 344546 115174
rect 344782 114938 344866 115174
rect 345102 114938 345134 115174
rect 344514 114854 345134 114938
rect 344514 114618 344546 114854
rect 344782 114618 344866 114854
rect 345102 114618 345134 114854
rect 344514 79174 345134 114618
rect 344514 78938 344546 79174
rect 344782 78938 344866 79174
rect 345102 78938 345134 79174
rect 344514 78854 345134 78938
rect 344514 78618 344546 78854
rect 344782 78618 344866 78854
rect 345102 78618 345134 78854
rect 344514 43174 345134 78618
rect 344514 42938 344546 43174
rect 344782 42938 344866 43174
rect 345102 42938 345134 43174
rect 344514 42854 345134 42938
rect 344514 42618 344546 42854
rect 344782 42618 344866 42854
rect 345102 42618 345134 42854
rect 344514 7174 345134 42618
rect 344514 6938 344546 7174
rect 344782 6938 344866 7174
rect 345102 6938 345134 7174
rect 344514 6854 345134 6938
rect 344514 6618 344546 6854
rect 344782 6618 344866 6854
rect 345102 6618 345134 6854
rect 344514 -2266 345134 6618
rect 344514 -2502 344546 -2266
rect 344782 -2502 344866 -2266
rect 345102 -2502 345134 -2266
rect 344514 -2586 345134 -2502
rect 344514 -2822 344546 -2586
rect 344782 -2822 344866 -2586
rect 345102 -2822 345134 -2586
rect 344514 -3814 345134 -2822
rect 348234 694894 348854 708122
rect 348234 694658 348266 694894
rect 348502 694658 348586 694894
rect 348822 694658 348854 694894
rect 348234 694574 348854 694658
rect 348234 694338 348266 694574
rect 348502 694338 348586 694574
rect 348822 694338 348854 694574
rect 348234 658894 348854 694338
rect 348234 658658 348266 658894
rect 348502 658658 348586 658894
rect 348822 658658 348854 658894
rect 348234 658574 348854 658658
rect 348234 658338 348266 658574
rect 348502 658338 348586 658574
rect 348822 658338 348854 658574
rect 348234 622894 348854 658338
rect 348234 622658 348266 622894
rect 348502 622658 348586 622894
rect 348822 622658 348854 622894
rect 348234 622574 348854 622658
rect 348234 622338 348266 622574
rect 348502 622338 348586 622574
rect 348822 622338 348854 622574
rect 348234 586894 348854 622338
rect 348234 586658 348266 586894
rect 348502 586658 348586 586894
rect 348822 586658 348854 586894
rect 348234 586574 348854 586658
rect 348234 586338 348266 586574
rect 348502 586338 348586 586574
rect 348822 586338 348854 586574
rect 348234 550894 348854 586338
rect 348234 550658 348266 550894
rect 348502 550658 348586 550894
rect 348822 550658 348854 550894
rect 348234 550574 348854 550658
rect 348234 550338 348266 550574
rect 348502 550338 348586 550574
rect 348822 550338 348854 550574
rect 348234 514894 348854 550338
rect 348234 514658 348266 514894
rect 348502 514658 348586 514894
rect 348822 514658 348854 514894
rect 348234 514574 348854 514658
rect 348234 514338 348266 514574
rect 348502 514338 348586 514574
rect 348822 514338 348854 514574
rect 348234 478894 348854 514338
rect 348234 478658 348266 478894
rect 348502 478658 348586 478894
rect 348822 478658 348854 478894
rect 348234 478574 348854 478658
rect 348234 478338 348266 478574
rect 348502 478338 348586 478574
rect 348822 478338 348854 478574
rect 348234 442894 348854 478338
rect 348234 442658 348266 442894
rect 348502 442658 348586 442894
rect 348822 442658 348854 442894
rect 348234 442574 348854 442658
rect 348234 442338 348266 442574
rect 348502 442338 348586 442574
rect 348822 442338 348854 442574
rect 348234 406894 348854 442338
rect 348234 406658 348266 406894
rect 348502 406658 348586 406894
rect 348822 406658 348854 406894
rect 348234 406574 348854 406658
rect 348234 406338 348266 406574
rect 348502 406338 348586 406574
rect 348822 406338 348854 406574
rect 348234 370894 348854 406338
rect 348234 370658 348266 370894
rect 348502 370658 348586 370894
rect 348822 370658 348854 370894
rect 348234 370574 348854 370658
rect 348234 370338 348266 370574
rect 348502 370338 348586 370574
rect 348822 370338 348854 370574
rect 348234 334894 348854 370338
rect 348234 334658 348266 334894
rect 348502 334658 348586 334894
rect 348822 334658 348854 334894
rect 348234 334574 348854 334658
rect 348234 334338 348266 334574
rect 348502 334338 348586 334574
rect 348822 334338 348854 334574
rect 348234 298894 348854 334338
rect 348234 298658 348266 298894
rect 348502 298658 348586 298894
rect 348822 298658 348854 298894
rect 348234 298574 348854 298658
rect 348234 298338 348266 298574
rect 348502 298338 348586 298574
rect 348822 298338 348854 298574
rect 348234 262894 348854 298338
rect 348234 262658 348266 262894
rect 348502 262658 348586 262894
rect 348822 262658 348854 262894
rect 348234 262574 348854 262658
rect 348234 262338 348266 262574
rect 348502 262338 348586 262574
rect 348822 262338 348854 262574
rect 348234 226894 348854 262338
rect 348234 226658 348266 226894
rect 348502 226658 348586 226894
rect 348822 226658 348854 226894
rect 348234 226574 348854 226658
rect 348234 226338 348266 226574
rect 348502 226338 348586 226574
rect 348822 226338 348854 226574
rect 348234 190894 348854 226338
rect 348234 190658 348266 190894
rect 348502 190658 348586 190894
rect 348822 190658 348854 190894
rect 348234 190574 348854 190658
rect 348234 190338 348266 190574
rect 348502 190338 348586 190574
rect 348822 190338 348854 190574
rect 348234 154894 348854 190338
rect 348234 154658 348266 154894
rect 348502 154658 348586 154894
rect 348822 154658 348854 154894
rect 348234 154574 348854 154658
rect 348234 154338 348266 154574
rect 348502 154338 348586 154574
rect 348822 154338 348854 154574
rect 348234 118894 348854 154338
rect 348234 118658 348266 118894
rect 348502 118658 348586 118894
rect 348822 118658 348854 118894
rect 348234 118574 348854 118658
rect 348234 118338 348266 118574
rect 348502 118338 348586 118574
rect 348822 118338 348854 118574
rect 348234 82894 348854 118338
rect 348234 82658 348266 82894
rect 348502 82658 348586 82894
rect 348822 82658 348854 82894
rect 348234 82574 348854 82658
rect 348234 82338 348266 82574
rect 348502 82338 348586 82574
rect 348822 82338 348854 82574
rect 348234 46894 348854 82338
rect 348234 46658 348266 46894
rect 348502 46658 348586 46894
rect 348822 46658 348854 46894
rect 348234 46574 348854 46658
rect 348234 46338 348266 46574
rect 348502 46338 348586 46574
rect 348822 46338 348854 46574
rect 348234 10894 348854 46338
rect 348234 10658 348266 10894
rect 348502 10658 348586 10894
rect 348822 10658 348854 10894
rect 348234 10574 348854 10658
rect 348234 10338 348266 10574
rect 348502 10338 348586 10574
rect 348822 10338 348854 10574
rect 348234 -4186 348854 10338
rect 350794 705798 351414 705830
rect 350794 705562 350826 705798
rect 351062 705562 351146 705798
rect 351382 705562 351414 705798
rect 350794 705478 351414 705562
rect 350794 705242 350826 705478
rect 351062 705242 351146 705478
rect 351382 705242 351414 705478
rect 350794 669454 351414 705242
rect 350794 669218 350826 669454
rect 351062 669218 351146 669454
rect 351382 669218 351414 669454
rect 350794 669134 351414 669218
rect 350794 668898 350826 669134
rect 351062 668898 351146 669134
rect 351382 668898 351414 669134
rect 350794 633454 351414 668898
rect 350794 633218 350826 633454
rect 351062 633218 351146 633454
rect 351382 633218 351414 633454
rect 350794 633134 351414 633218
rect 350794 632898 350826 633134
rect 351062 632898 351146 633134
rect 351382 632898 351414 633134
rect 350794 597454 351414 632898
rect 350794 597218 350826 597454
rect 351062 597218 351146 597454
rect 351382 597218 351414 597454
rect 350794 597134 351414 597218
rect 350794 596898 350826 597134
rect 351062 596898 351146 597134
rect 351382 596898 351414 597134
rect 350794 561454 351414 596898
rect 350794 561218 350826 561454
rect 351062 561218 351146 561454
rect 351382 561218 351414 561454
rect 350794 561134 351414 561218
rect 350794 560898 350826 561134
rect 351062 560898 351146 561134
rect 351382 560898 351414 561134
rect 350794 525454 351414 560898
rect 350794 525218 350826 525454
rect 351062 525218 351146 525454
rect 351382 525218 351414 525454
rect 350794 525134 351414 525218
rect 350794 524898 350826 525134
rect 351062 524898 351146 525134
rect 351382 524898 351414 525134
rect 350794 489454 351414 524898
rect 350794 489218 350826 489454
rect 351062 489218 351146 489454
rect 351382 489218 351414 489454
rect 350794 489134 351414 489218
rect 350794 488898 350826 489134
rect 351062 488898 351146 489134
rect 351382 488898 351414 489134
rect 350794 453454 351414 488898
rect 350794 453218 350826 453454
rect 351062 453218 351146 453454
rect 351382 453218 351414 453454
rect 350794 453134 351414 453218
rect 350794 452898 350826 453134
rect 351062 452898 351146 453134
rect 351382 452898 351414 453134
rect 350794 417454 351414 452898
rect 350794 417218 350826 417454
rect 351062 417218 351146 417454
rect 351382 417218 351414 417454
rect 350794 417134 351414 417218
rect 350794 416898 350826 417134
rect 351062 416898 351146 417134
rect 351382 416898 351414 417134
rect 350794 381454 351414 416898
rect 350794 381218 350826 381454
rect 351062 381218 351146 381454
rect 351382 381218 351414 381454
rect 350794 381134 351414 381218
rect 350794 380898 350826 381134
rect 351062 380898 351146 381134
rect 351382 380898 351414 381134
rect 350794 345454 351414 380898
rect 350794 345218 350826 345454
rect 351062 345218 351146 345454
rect 351382 345218 351414 345454
rect 350794 345134 351414 345218
rect 350794 344898 350826 345134
rect 351062 344898 351146 345134
rect 351382 344898 351414 345134
rect 350794 309454 351414 344898
rect 350794 309218 350826 309454
rect 351062 309218 351146 309454
rect 351382 309218 351414 309454
rect 350794 309134 351414 309218
rect 350794 308898 350826 309134
rect 351062 308898 351146 309134
rect 351382 308898 351414 309134
rect 350794 273454 351414 308898
rect 350794 273218 350826 273454
rect 351062 273218 351146 273454
rect 351382 273218 351414 273454
rect 350794 273134 351414 273218
rect 350794 272898 350826 273134
rect 351062 272898 351146 273134
rect 351382 272898 351414 273134
rect 350794 237454 351414 272898
rect 350794 237218 350826 237454
rect 351062 237218 351146 237454
rect 351382 237218 351414 237454
rect 350794 237134 351414 237218
rect 350794 236898 350826 237134
rect 351062 236898 351146 237134
rect 351382 236898 351414 237134
rect 350794 201454 351414 236898
rect 350794 201218 350826 201454
rect 351062 201218 351146 201454
rect 351382 201218 351414 201454
rect 350794 201134 351414 201218
rect 350794 200898 350826 201134
rect 351062 200898 351146 201134
rect 351382 200898 351414 201134
rect 350794 165454 351414 200898
rect 350794 165218 350826 165454
rect 351062 165218 351146 165454
rect 351382 165218 351414 165454
rect 350794 165134 351414 165218
rect 350794 164898 350826 165134
rect 351062 164898 351146 165134
rect 351382 164898 351414 165134
rect 350794 129454 351414 164898
rect 350794 129218 350826 129454
rect 351062 129218 351146 129454
rect 351382 129218 351414 129454
rect 350794 129134 351414 129218
rect 350794 128898 350826 129134
rect 351062 128898 351146 129134
rect 351382 128898 351414 129134
rect 350794 93454 351414 128898
rect 350794 93218 350826 93454
rect 351062 93218 351146 93454
rect 351382 93218 351414 93454
rect 350794 93134 351414 93218
rect 350794 92898 350826 93134
rect 351062 92898 351146 93134
rect 351382 92898 351414 93134
rect 350794 57454 351414 92898
rect 350794 57218 350826 57454
rect 351062 57218 351146 57454
rect 351382 57218 351414 57454
rect 350794 57134 351414 57218
rect 350794 56898 350826 57134
rect 351062 56898 351146 57134
rect 351382 56898 351414 57134
rect 350794 21454 351414 56898
rect 350794 21218 350826 21454
rect 351062 21218 351146 21454
rect 351382 21218 351414 21454
rect 350794 21134 351414 21218
rect 350794 20898 350826 21134
rect 351062 20898 351146 21134
rect 351382 20898 351414 21134
rect 350794 -1306 351414 20898
rect 350794 -1542 350826 -1306
rect 351062 -1542 351146 -1306
rect 351382 -1542 351414 -1306
rect 350794 -1626 351414 -1542
rect 350794 -1862 350826 -1626
rect 351062 -1862 351146 -1626
rect 351382 -1862 351414 -1626
rect 350794 -1894 351414 -1862
rect 351954 698614 352574 710042
rect 361954 711558 362574 711590
rect 361954 711322 361986 711558
rect 362222 711322 362306 711558
rect 362542 711322 362574 711558
rect 361954 711238 362574 711322
rect 361954 711002 361986 711238
rect 362222 711002 362306 711238
rect 362542 711002 362574 711238
rect 358234 709638 358854 709670
rect 358234 709402 358266 709638
rect 358502 709402 358586 709638
rect 358822 709402 358854 709638
rect 358234 709318 358854 709402
rect 358234 709082 358266 709318
rect 358502 709082 358586 709318
rect 358822 709082 358854 709318
rect 351954 698378 351986 698614
rect 352222 698378 352306 698614
rect 352542 698378 352574 698614
rect 351954 698294 352574 698378
rect 351954 698058 351986 698294
rect 352222 698058 352306 698294
rect 352542 698058 352574 698294
rect 351954 662614 352574 698058
rect 351954 662378 351986 662614
rect 352222 662378 352306 662614
rect 352542 662378 352574 662614
rect 351954 662294 352574 662378
rect 351954 662058 351986 662294
rect 352222 662058 352306 662294
rect 352542 662058 352574 662294
rect 351954 626614 352574 662058
rect 351954 626378 351986 626614
rect 352222 626378 352306 626614
rect 352542 626378 352574 626614
rect 351954 626294 352574 626378
rect 351954 626058 351986 626294
rect 352222 626058 352306 626294
rect 352542 626058 352574 626294
rect 351954 590614 352574 626058
rect 351954 590378 351986 590614
rect 352222 590378 352306 590614
rect 352542 590378 352574 590614
rect 351954 590294 352574 590378
rect 351954 590058 351986 590294
rect 352222 590058 352306 590294
rect 352542 590058 352574 590294
rect 351954 554614 352574 590058
rect 351954 554378 351986 554614
rect 352222 554378 352306 554614
rect 352542 554378 352574 554614
rect 351954 554294 352574 554378
rect 351954 554058 351986 554294
rect 352222 554058 352306 554294
rect 352542 554058 352574 554294
rect 351954 518614 352574 554058
rect 351954 518378 351986 518614
rect 352222 518378 352306 518614
rect 352542 518378 352574 518614
rect 351954 518294 352574 518378
rect 351954 518058 351986 518294
rect 352222 518058 352306 518294
rect 352542 518058 352574 518294
rect 351954 482614 352574 518058
rect 351954 482378 351986 482614
rect 352222 482378 352306 482614
rect 352542 482378 352574 482614
rect 351954 482294 352574 482378
rect 351954 482058 351986 482294
rect 352222 482058 352306 482294
rect 352542 482058 352574 482294
rect 351954 446614 352574 482058
rect 351954 446378 351986 446614
rect 352222 446378 352306 446614
rect 352542 446378 352574 446614
rect 351954 446294 352574 446378
rect 351954 446058 351986 446294
rect 352222 446058 352306 446294
rect 352542 446058 352574 446294
rect 351954 410614 352574 446058
rect 351954 410378 351986 410614
rect 352222 410378 352306 410614
rect 352542 410378 352574 410614
rect 351954 410294 352574 410378
rect 351954 410058 351986 410294
rect 352222 410058 352306 410294
rect 352542 410058 352574 410294
rect 351954 374614 352574 410058
rect 351954 374378 351986 374614
rect 352222 374378 352306 374614
rect 352542 374378 352574 374614
rect 351954 374294 352574 374378
rect 351954 374058 351986 374294
rect 352222 374058 352306 374294
rect 352542 374058 352574 374294
rect 351954 338614 352574 374058
rect 351954 338378 351986 338614
rect 352222 338378 352306 338614
rect 352542 338378 352574 338614
rect 351954 338294 352574 338378
rect 351954 338058 351986 338294
rect 352222 338058 352306 338294
rect 352542 338058 352574 338294
rect 351954 302614 352574 338058
rect 351954 302378 351986 302614
rect 352222 302378 352306 302614
rect 352542 302378 352574 302614
rect 351954 302294 352574 302378
rect 351954 302058 351986 302294
rect 352222 302058 352306 302294
rect 352542 302058 352574 302294
rect 351954 266614 352574 302058
rect 351954 266378 351986 266614
rect 352222 266378 352306 266614
rect 352542 266378 352574 266614
rect 351954 266294 352574 266378
rect 351954 266058 351986 266294
rect 352222 266058 352306 266294
rect 352542 266058 352574 266294
rect 351954 230614 352574 266058
rect 351954 230378 351986 230614
rect 352222 230378 352306 230614
rect 352542 230378 352574 230614
rect 351954 230294 352574 230378
rect 351954 230058 351986 230294
rect 352222 230058 352306 230294
rect 352542 230058 352574 230294
rect 351954 194614 352574 230058
rect 351954 194378 351986 194614
rect 352222 194378 352306 194614
rect 352542 194378 352574 194614
rect 351954 194294 352574 194378
rect 351954 194058 351986 194294
rect 352222 194058 352306 194294
rect 352542 194058 352574 194294
rect 351954 158614 352574 194058
rect 351954 158378 351986 158614
rect 352222 158378 352306 158614
rect 352542 158378 352574 158614
rect 351954 158294 352574 158378
rect 351954 158058 351986 158294
rect 352222 158058 352306 158294
rect 352542 158058 352574 158294
rect 351954 122614 352574 158058
rect 351954 122378 351986 122614
rect 352222 122378 352306 122614
rect 352542 122378 352574 122614
rect 351954 122294 352574 122378
rect 351954 122058 351986 122294
rect 352222 122058 352306 122294
rect 352542 122058 352574 122294
rect 351954 86614 352574 122058
rect 351954 86378 351986 86614
rect 352222 86378 352306 86614
rect 352542 86378 352574 86614
rect 351954 86294 352574 86378
rect 351954 86058 351986 86294
rect 352222 86058 352306 86294
rect 352542 86058 352574 86294
rect 351954 50614 352574 86058
rect 351954 50378 351986 50614
rect 352222 50378 352306 50614
rect 352542 50378 352574 50614
rect 351954 50294 352574 50378
rect 351954 50058 351986 50294
rect 352222 50058 352306 50294
rect 352542 50058 352574 50294
rect 351954 14614 352574 50058
rect 351954 14378 351986 14614
rect 352222 14378 352306 14614
rect 352542 14378 352574 14614
rect 351954 14294 352574 14378
rect 351954 14058 351986 14294
rect 352222 14058 352306 14294
rect 352542 14058 352574 14294
rect 348234 -4422 348266 -4186
rect 348502 -4422 348586 -4186
rect 348822 -4422 348854 -4186
rect 348234 -4506 348854 -4422
rect 348234 -4742 348266 -4506
rect 348502 -4742 348586 -4506
rect 348822 -4742 348854 -4506
rect 348234 -5734 348854 -4742
rect 341954 -7302 341986 -7066
rect 342222 -7302 342306 -7066
rect 342542 -7302 342574 -7066
rect 341954 -7386 342574 -7302
rect 341954 -7622 341986 -7386
rect 342222 -7622 342306 -7386
rect 342542 -7622 342574 -7386
rect 341954 -7654 342574 -7622
rect 351954 -6106 352574 14058
rect 354514 707718 355134 707750
rect 354514 707482 354546 707718
rect 354782 707482 354866 707718
rect 355102 707482 355134 707718
rect 354514 707398 355134 707482
rect 354514 707162 354546 707398
rect 354782 707162 354866 707398
rect 355102 707162 355134 707398
rect 354514 673174 355134 707162
rect 354514 672938 354546 673174
rect 354782 672938 354866 673174
rect 355102 672938 355134 673174
rect 354514 672854 355134 672938
rect 354514 672618 354546 672854
rect 354782 672618 354866 672854
rect 355102 672618 355134 672854
rect 354514 637174 355134 672618
rect 354514 636938 354546 637174
rect 354782 636938 354866 637174
rect 355102 636938 355134 637174
rect 354514 636854 355134 636938
rect 354514 636618 354546 636854
rect 354782 636618 354866 636854
rect 355102 636618 355134 636854
rect 354514 601174 355134 636618
rect 354514 600938 354546 601174
rect 354782 600938 354866 601174
rect 355102 600938 355134 601174
rect 354514 600854 355134 600938
rect 354514 600618 354546 600854
rect 354782 600618 354866 600854
rect 355102 600618 355134 600854
rect 354514 565174 355134 600618
rect 354514 564938 354546 565174
rect 354782 564938 354866 565174
rect 355102 564938 355134 565174
rect 354514 564854 355134 564938
rect 354514 564618 354546 564854
rect 354782 564618 354866 564854
rect 355102 564618 355134 564854
rect 354514 529174 355134 564618
rect 354514 528938 354546 529174
rect 354782 528938 354866 529174
rect 355102 528938 355134 529174
rect 354514 528854 355134 528938
rect 354514 528618 354546 528854
rect 354782 528618 354866 528854
rect 355102 528618 355134 528854
rect 354514 493174 355134 528618
rect 354514 492938 354546 493174
rect 354782 492938 354866 493174
rect 355102 492938 355134 493174
rect 354514 492854 355134 492938
rect 354514 492618 354546 492854
rect 354782 492618 354866 492854
rect 355102 492618 355134 492854
rect 354514 457174 355134 492618
rect 354514 456938 354546 457174
rect 354782 456938 354866 457174
rect 355102 456938 355134 457174
rect 354514 456854 355134 456938
rect 354514 456618 354546 456854
rect 354782 456618 354866 456854
rect 355102 456618 355134 456854
rect 354514 421174 355134 456618
rect 354514 420938 354546 421174
rect 354782 420938 354866 421174
rect 355102 420938 355134 421174
rect 354514 420854 355134 420938
rect 354514 420618 354546 420854
rect 354782 420618 354866 420854
rect 355102 420618 355134 420854
rect 354514 385174 355134 420618
rect 354514 384938 354546 385174
rect 354782 384938 354866 385174
rect 355102 384938 355134 385174
rect 354514 384854 355134 384938
rect 354514 384618 354546 384854
rect 354782 384618 354866 384854
rect 355102 384618 355134 384854
rect 354514 349174 355134 384618
rect 354514 348938 354546 349174
rect 354782 348938 354866 349174
rect 355102 348938 355134 349174
rect 354514 348854 355134 348938
rect 354514 348618 354546 348854
rect 354782 348618 354866 348854
rect 355102 348618 355134 348854
rect 354514 313174 355134 348618
rect 354514 312938 354546 313174
rect 354782 312938 354866 313174
rect 355102 312938 355134 313174
rect 354514 312854 355134 312938
rect 354514 312618 354546 312854
rect 354782 312618 354866 312854
rect 355102 312618 355134 312854
rect 354514 277174 355134 312618
rect 354514 276938 354546 277174
rect 354782 276938 354866 277174
rect 355102 276938 355134 277174
rect 354514 276854 355134 276938
rect 354514 276618 354546 276854
rect 354782 276618 354866 276854
rect 355102 276618 355134 276854
rect 354514 241174 355134 276618
rect 354514 240938 354546 241174
rect 354782 240938 354866 241174
rect 355102 240938 355134 241174
rect 354514 240854 355134 240938
rect 354514 240618 354546 240854
rect 354782 240618 354866 240854
rect 355102 240618 355134 240854
rect 354514 205174 355134 240618
rect 354514 204938 354546 205174
rect 354782 204938 354866 205174
rect 355102 204938 355134 205174
rect 354514 204854 355134 204938
rect 354514 204618 354546 204854
rect 354782 204618 354866 204854
rect 355102 204618 355134 204854
rect 354514 169174 355134 204618
rect 354514 168938 354546 169174
rect 354782 168938 354866 169174
rect 355102 168938 355134 169174
rect 354514 168854 355134 168938
rect 354514 168618 354546 168854
rect 354782 168618 354866 168854
rect 355102 168618 355134 168854
rect 354514 133174 355134 168618
rect 354514 132938 354546 133174
rect 354782 132938 354866 133174
rect 355102 132938 355134 133174
rect 354514 132854 355134 132938
rect 354514 132618 354546 132854
rect 354782 132618 354866 132854
rect 355102 132618 355134 132854
rect 354514 97174 355134 132618
rect 354514 96938 354546 97174
rect 354782 96938 354866 97174
rect 355102 96938 355134 97174
rect 354514 96854 355134 96938
rect 354514 96618 354546 96854
rect 354782 96618 354866 96854
rect 355102 96618 355134 96854
rect 354514 61174 355134 96618
rect 354514 60938 354546 61174
rect 354782 60938 354866 61174
rect 355102 60938 355134 61174
rect 354514 60854 355134 60938
rect 354514 60618 354546 60854
rect 354782 60618 354866 60854
rect 355102 60618 355134 60854
rect 354514 25174 355134 60618
rect 354514 24938 354546 25174
rect 354782 24938 354866 25174
rect 355102 24938 355134 25174
rect 354514 24854 355134 24938
rect 354514 24618 354546 24854
rect 354782 24618 354866 24854
rect 355102 24618 355134 24854
rect 354514 -3226 355134 24618
rect 354514 -3462 354546 -3226
rect 354782 -3462 354866 -3226
rect 355102 -3462 355134 -3226
rect 354514 -3546 355134 -3462
rect 354514 -3782 354546 -3546
rect 354782 -3782 354866 -3546
rect 355102 -3782 355134 -3546
rect 354514 -3814 355134 -3782
rect 358234 676894 358854 709082
rect 358234 676658 358266 676894
rect 358502 676658 358586 676894
rect 358822 676658 358854 676894
rect 358234 676574 358854 676658
rect 358234 676338 358266 676574
rect 358502 676338 358586 676574
rect 358822 676338 358854 676574
rect 358234 640894 358854 676338
rect 358234 640658 358266 640894
rect 358502 640658 358586 640894
rect 358822 640658 358854 640894
rect 358234 640574 358854 640658
rect 358234 640338 358266 640574
rect 358502 640338 358586 640574
rect 358822 640338 358854 640574
rect 358234 604894 358854 640338
rect 358234 604658 358266 604894
rect 358502 604658 358586 604894
rect 358822 604658 358854 604894
rect 358234 604574 358854 604658
rect 358234 604338 358266 604574
rect 358502 604338 358586 604574
rect 358822 604338 358854 604574
rect 358234 568894 358854 604338
rect 358234 568658 358266 568894
rect 358502 568658 358586 568894
rect 358822 568658 358854 568894
rect 358234 568574 358854 568658
rect 358234 568338 358266 568574
rect 358502 568338 358586 568574
rect 358822 568338 358854 568574
rect 358234 532894 358854 568338
rect 358234 532658 358266 532894
rect 358502 532658 358586 532894
rect 358822 532658 358854 532894
rect 358234 532574 358854 532658
rect 358234 532338 358266 532574
rect 358502 532338 358586 532574
rect 358822 532338 358854 532574
rect 358234 496894 358854 532338
rect 358234 496658 358266 496894
rect 358502 496658 358586 496894
rect 358822 496658 358854 496894
rect 358234 496574 358854 496658
rect 358234 496338 358266 496574
rect 358502 496338 358586 496574
rect 358822 496338 358854 496574
rect 358234 460894 358854 496338
rect 358234 460658 358266 460894
rect 358502 460658 358586 460894
rect 358822 460658 358854 460894
rect 358234 460574 358854 460658
rect 358234 460338 358266 460574
rect 358502 460338 358586 460574
rect 358822 460338 358854 460574
rect 358234 424894 358854 460338
rect 358234 424658 358266 424894
rect 358502 424658 358586 424894
rect 358822 424658 358854 424894
rect 358234 424574 358854 424658
rect 358234 424338 358266 424574
rect 358502 424338 358586 424574
rect 358822 424338 358854 424574
rect 358234 388894 358854 424338
rect 358234 388658 358266 388894
rect 358502 388658 358586 388894
rect 358822 388658 358854 388894
rect 358234 388574 358854 388658
rect 358234 388338 358266 388574
rect 358502 388338 358586 388574
rect 358822 388338 358854 388574
rect 358234 352894 358854 388338
rect 358234 352658 358266 352894
rect 358502 352658 358586 352894
rect 358822 352658 358854 352894
rect 358234 352574 358854 352658
rect 358234 352338 358266 352574
rect 358502 352338 358586 352574
rect 358822 352338 358854 352574
rect 358234 316894 358854 352338
rect 358234 316658 358266 316894
rect 358502 316658 358586 316894
rect 358822 316658 358854 316894
rect 358234 316574 358854 316658
rect 358234 316338 358266 316574
rect 358502 316338 358586 316574
rect 358822 316338 358854 316574
rect 358234 280894 358854 316338
rect 358234 280658 358266 280894
rect 358502 280658 358586 280894
rect 358822 280658 358854 280894
rect 358234 280574 358854 280658
rect 358234 280338 358266 280574
rect 358502 280338 358586 280574
rect 358822 280338 358854 280574
rect 358234 244894 358854 280338
rect 358234 244658 358266 244894
rect 358502 244658 358586 244894
rect 358822 244658 358854 244894
rect 358234 244574 358854 244658
rect 358234 244338 358266 244574
rect 358502 244338 358586 244574
rect 358822 244338 358854 244574
rect 358234 208894 358854 244338
rect 358234 208658 358266 208894
rect 358502 208658 358586 208894
rect 358822 208658 358854 208894
rect 358234 208574 358854 208658
rect 358234 208338 358266 208574
rect 358502 208338 358586 208574
rect 358822 208338 358854 208574
rect 358234 172894 358854 208338
rect 358234 172658 358266 172894
rect 358502 172658 358586 172894
rect 358822 172658 358854 172894
rect 358234 172574 358854 172658
rect 358234 172338 358266 172574
rect 358502 172338 358586 172574
rect 358822 172338 358854 172574
rect 358234 136894 358854 172338
rect 358234 136658 358266 136894
rect 358502 136658 358586 136894
rect 358822 136658 358854 136894
rect 358234 136574 358854 136658
rect 358234 136338 358266 136574
rect 358502 136338 358586 136574
rect 358822 136338 358854 136574
rect 358234 100894 358854 136338
rect 358234 100658 358266 100894
rect 358502 100658 358586 100894
rect 358822 100658 358854 100894
rect 358234 100574 358854 100658
rect 358234 100338 358266 100574
rect 358502 100338 358586 100574
rect 358822 100338 358854 100574
rect 358234 64894 358854 100338
rect 358234 64658 358266 64894
rect 358502 64658 358586 64894
rect 358822 64658 358854 64894
rect 358234 64574 358854 64658
rect 358234 64338 358266 64574
rect 358502 64338 358586 64574
rect 358822 64338 358854 64574
rect 358234 28894 358854 64338
rect 358234 28658 358266 28894
rect 358502 28658 358586 28894
rect 358822 28658 358854 28894
rect 358234 28574 358854 28658
rect 358234 28338 358266 28574
rect 358502 28338 358586 28574
rect 358822 28338 358854 28574
rect 358234 -5146 358854 28338
rect 360794 704838 361414 705830
rect 360794 704602 360826 704838
rect 361062 704602 361146 704838
rect 361382 704602 361414 704838
rect 360794 704518 361414 704602
rect 360794 704282 360826 704518
rect 361062 704282 361146 704518
rect 361382 704282 361414 704518
rect 360794 687454 361414 704282
rect 360794 687218 360826 687454
rect 361062 687218 361146 687454
rect 361382 687218 361414 687454
rect 360794 687134 361414 687218
rect 360794 686898 360826 687134
rect 361062 686898 361146 687134
rect 361382 686898 361414 687134
rect 360794 651454 361414 686898
rect 360794 651218 360826 651454
rect 361062 651218 361146 651454
rect 361382 651218 361414 651454
rect 360794 651134 361414 651218
rect 360794 650898 360826 651134
rect 361062 650898 361146 651134
rect 361382 650898 361414 651134
rect 360794 615454 361414 650898
rect 360794 615218 360826 615454
rect 361062 615218 361146 615454
rect 361382 615218 361414 615454
rect 360794 615134 361414 615218
rect 360794 614898 360826 615134
rect 361062 614898 361146 615134
rect 361382 614898 361414 615134
rect 360794 579454 361414 614898
rect 360794 579218 360826 579454
rect 361062 579218 361146 579454
rect 361382 579218 361414 579454
rect 360794 579134 361414 579218
rect 360794 578898 360826 579134
rect 361062 578898 361146 579134
rect 361382 578898 361414 579134
rect 360794 543454 361414 578898
rect 360794 543218 360826 543454
rect 361062 543218 361146 543454
rect 361382 543218 361414 543454
rect 360794 543134 361414 543218
rect 360794 542898 360826 543134
rect 361062 542898 361146 543134
rect 361382 542898 361414 543134
rect 360794 507454 361414 542898
rect 360794 507218 360826 507454
rect 361062 507218 361146 507454
rect 361382 507218 361414 507454
rect 360794 507134 361414 507218
rect 360794 506898 360826 507134
rect 361062 506898 361146 507134
rect 361382 506898 361414 507134
rect 360794 471454 361414 506898
rect 360794 471218 360826 471454
rect 361062 471218 361146 471454
rect 361382 471218 361414 471454
rect 360794 471134 361414 471218
rect 360794 470898 360826 471134
rect 361062 470898 361146 471134
rect 361382 470898 361414 471134
rect 360794 435454 361414 470898
rect 360794 435218 360826 435454
rect 361062 435218 361146 435454
rect 361382 435218 361414 435454
rect 360794 435134 361414 435218
rect 360794 434898 360826 435134
rect 361062 434898 361146 435134
rect 361382 434898 361414 435134
rect 360794 399454 361414 434898
rect 360794 399218 360826 399454
rect 361062 399218 361146 399454
rect 361382 399218 361414 399454
rect 360794 399134 361414 399218
rect 360794 398898 360826 399134
rect 361062 398898 361146 399134
rect 361382 398898 361414 399134
rect 360794 363454 361414 398898
rect 360794 363218 360826 363454
rect 361062 363218 361146 363454
rect 361382 363218 361414 363454
rect 360794 363134 361414 363218
rect 360794 362898 360826 363134
rect 361062 362898 361146 363134
rect 361382 362898 361414 363134
rect 360794 327454 361414 362898
rect 360794 327218 360826 327454
rect 361062 327218 361146 327454
rect 361382 327218 361414 327454
rect 360794 327134 361414 327218
rect 360794 326898 360826 327134
rect 361062 326898 361146 327134
rect 361382 326898 361414 327134
rect 360794 291454 361414 326898
rect 360794 291218 360826 291454
rect 361062 291218 361146 291454
rect 361382 291218 361414 291454
rect 360794 291134 361414 291218
rect 360794 290898 360826 291134
rect 361062 290898 361146 291134
rect 361382 290898 361414 291134
rect 360794 255454 361414 290898
rect 360794 255218 360826 255454
rect 361062 255218 361146 255454
rect 361382 255218 361414 255454
rect 360794 255134 361414 255218
rect 360794 254898 360826 255134
rect 361062 254898 361146 255134
rect 361382 254898 361414 255134
rect 360794 219454 361414 254898
rect 360794 219218 360826 219454
rect 361062 219218 361146 219454
rect 361382 219218 361414 219454
rect 360794 219134 361414 219218
rect 360794 218898 360826 219134
rect 361062 218898 361146 219134
rect 361382 218898 361414 219134
rect 360794 183454 361414 218898
rect 360794 183218 360826 183454
rect 361062 183218 361146 183454
rect 361382 183218 361414 183454
rect 360794 183134 361414 183218
rect 360794 182898 360826 183134
rect 361062 182898 361146 183134
rect 361382 182898 361414 183134
rect 360794 147454 361414 182898
rect 360794 147218 360826 147454
rect 361062 147218 361146 147454
rect 361382 147218 361414 147454
rect 360794 147134 361414 147218
rect 360794 146898 360826 147134
rect 361062 146898 361146 147134
rect 361382 146898 361414 147134
rect 360794 111454 361414 146898
rect 360794 111218 360826 111454
rect 361062 111218 361146 111454
rect 361382 111218 361414 111454
rect 360794 111134 361414 111218
rect 360794 110898 360826 111134
rect 361062 110898 361146 111134
rect 361382 110898 361414 111134
rect 360794 75454 361414 110898
rect 360794 75218 360826 75454
rect 361062 75218 361146 75454
rect 361382 75218 361414 75454
rect 360794 75134 361414 75218
rect 360794 74898 360826 75134
rect 361062 74898 361146 75134
rect 361382 74898 361414 75134
rect 360794 39454 361414 74898
rect 360794 39218 360826 39454
rect 361062 39218 361146 39454
rect 361382 39218 361414 39454
rect 360794 39134 361414 39218
rect 360794 38898 360826 39134
rect 361062 38898 361146 39134
rect 361382 38898 361414 39134
rect 360794 3454 361414 38898
rect 360794 3218 360826 3454
rect 361062 3218 361146 3454
rect 361382 3218 361414 3454
rect 360794 3134 361414 3218
rect 360794 2898 360826 3134
rect 361062 2898 361146 3134
rect 361382 2898 361414 3134
rect 360794 -346 361414 2898
rect 360794 -582 360826 -346
rect 361062 -582 361146 -346
rect 361382 -582 361414 -346
rect 360794 -666 361414 -582
rect 360794 -902 360826 -666
rect 361062 -902 361146 -666
rect 361382 -902 361414 -666
rect 360794 -1894 361414 -902
rect 361954 680614 362574 711002
rect 371954 710598 372574 711590
rect 371954 710362 371986 710598
rect 372222 710362 372306 710598
rect 372542 710362 372574 710598
rect 371954 710278 372574 710362
rect 371954 710042 371986 710278
rect 372222 710042 372306 710278
rect 372542 710042 372574 710278
rect 368234 708678 368854 709670
rect 368234 708442 368266 708678
rect 368502 708442 368586 708678
rect 368822 708442 368854 708678
rect 368234 708358 368854 708442
rect 368234 708122 368266 708358
rect 368502 708122 368586 708358
rect 368822 708122 368854 708358
rect 361954 680378 361986 680614
rect 362222 680378 362306 680614
rect 362542 680378 362574 680614
rect 361954 680294 362574 680378
rect 361954 680058 361986 680294
rect 362222 680058 362306 680294
rect 362542 680058 362574 680294
rect 361954 644614 362574 680058
rect 361954 644378 361986 644614
rect 362222 644378 362306 644614
rect 362542 644378 362574 644614
rect 361954 644294 362574 644378
rect 361954 644058 361986 644294
rect 362222 644058 362306 644294
rect 362542 644058 362574 644294
rect 361954 608614 362574 644058
rect 361954 608378 361986 608614
rect 362222 608378 362306 608614
rect 362542 608378 362574 608614
rect 361954 608294 362574 608378
rect 361954 608058 361986 608294
rect 362222 608058 362306 608294
rect 362542 608058 362574 608294
rect 361954 572614 362574 608058
rect 361954 572378 361986 572614
rect 362222 572378 362306 572614
rect 362542 572378 362574 572614
rect 361954 572294 362574 572378
rect 361954 572058 361986 572294
rect 362222 572058 362306 572294
rect 362542 572058 362574 572294
rect 361954 536614 362574 572058
rect 361954 536378 361986 536614
rect 362222 536378 362306 536614
rect 362542 536378 362574 536614
rect 361954 536294 362574 536378
rect 361954 536058 361986 536294
rect 362222 536058 362306 536294
rect 362542 536058 362574 536294
rect 361954 500614 362574 536058
rect 361954 500378 361986 500614
rect 362222 500378 362306 500614
rect 362542 500378 362574 500614
rect 361954 500294 362574 500378
rect 361954 500058 361986 500294
rect 362222 500058 362306 500294
rect 362542 500058 362574 500294
rect 361954 464614 362574 500058
rect 361954 464378 361986 464614
rect 362222 464378 362306 464614
rect 362542 464378 362574 464614
rect 361954 464294 362574 464378
rect 361954 464058 361986 464294
rect 362222 464058 362306 464294
rect 362542 464058 362574 464294
rect 361954 428614 362574 464058
rect 361954 428378 361986 428614
rect 362222 428378 362306 428614
rect 362542 428378 362574 428614
rect 361954 428294 362574 428378
rect 361954 428058 361986 428294
rect 362222 428058 362306 428294
rect 362542 428058 362574 428294
rect 361954 392614 362574 428058
rect 361954 392378 361986 392614
rect 362222 392378 362306 392614
rect 362542 392378 362574 392614
rect 361954 392294 362574 392378
rect 361954 392058 361986 392294
rect 362222 392058 362306 392294
rect 362542 392058 362574 392294
rect 361954 356614 362574 392058
rect 361954 356378 361986 356614
rect 362222 356378 362306 356614
rect 362542 356378 362574 356614
rect 361954 356294 362574 356378
rect 361954 356058 361986 356294
rect 362222 356058 362306 356294
rect 362542 356058 362574 356294
rect 361954 320614 362574 356058
rect 361954 320378 361986 320614
rect 362222 320378 362306 320614
rect 362542 320378 362574 320614
rect 361954 320294 362574 320378
rect 361954 320058 361986 320294
rect 362222 320058 362306 320294
rect 362542 320058 362574 320294
rect 361954 284614 362574 320058
rect 361954 284378 361986 284614
rect 362222 284378 362306 284614
rect 362542 284378 362574 284614
rect 361954 284294 362574 284378
rect 361954 284058 361986 284294
rect 362222 284058 362306 284294
rect 362542 284058 362574 284294
rect 361954 248614 362574 284058
rect 361954 248378 361986 248614
rect 362222 248378 362306 248614
rect 362542 248378 362574 248614
rect 361954 248294 362574 248378
rect 361954 248058 361986 248294
rect 362222 248058 362306 248294
rect 362542 248058 362574 248294
rect 361954 212614 362574 248058
rect 361954 212378 361986 212614
rect 362222 212378 362306 212614
rect 362542 212378 362574 212614
rect 361954 212294 362574 212378
rect 361954 212058 361986 212294
rect 362222 212058 362306 212294
rect 362542 212058 362574 212294
rect 361954 176614 362574 212058
rect 361954 176378 361986 176614
rect 362222 176378 362306 176614
rect 362542 176378 362574 176614
rect 361954 176294 362574 176378
rect 361954 176058 361986 176294
rect 362222 176058 362306 176294
rect 362542 176058 362574 176294
rect 361954 140614 362574 176058
rect 361954 140378 361986 140614
rect 362222 140378 362306 140614
rect 362542 140378 362574 140614
rect 361954 140294 362574 140378
rect 361954 140058 361986 140294
rect 362222 140058 362306 140294
rect 362542 140058 362574 140294
rect 361954 104614 362574 140058
rect 361954 104378 361986 104614
rect 362222 104378 362306 104614
rect 362542 104378 362574 104614
rect 361954 104294 362574 104378
rect 361954 104058 361986 104294
rect 362222 104058 362306 104294
rect 362542 104058 362574 104294
rect 361954 68614 362574 104058
rect 361954 68378 361986 68614
rect 362222 68378 362306 68614
rect 362542 68378 362574 68614
rect 361954 68294 362574 68378
rect 361954 68058 361986 68294
rect 362222 68058 362306 68294
rect 362542 68058 362574 68294
rect 361954 32614 362574 68058
rect 361954 32378 361986 32614
rect 362222 32378 362306 32614
rect 362542 32378 362574 32614
rect 361954 32294 362574 32378
rect 361954 32058 361986 32294
rect 362222 32058 362306 32294
rect 362542 32058 362574 32294
rect 358234 -5382 358266 -5146
rect 358502 -5382 358586 -5146
rect 358822 -5382 358854 -5146
rect 358234 -5466 358854 -5382
rect 358234 -5702 358266 -5466
rect 358502 -5702 358586 -5466
rect 358822 -5702 358854 -5466
rect 358234 -5734 358854 -5702
rect 351954 -6342 351986 -6106
rect 352222 -6342 352306 -6106
rect 352542 -6342 352574 -6106
rect 351954 -6426 352574 -6342
rect 351954 -6662 351986 -6426
rect 352222 -6662 352306 -6426
rect 352542 -6662 352574 -6426
rect 351954 -7654 352574 -6662
rect 361954 -7066 362574 32058
rect 364514 706758 365134 707750
rect 364514 706522 364546 706758
rect 364782 706522 364866 706758
rect 365102 706522 365134 706758
rect 364514 706438 365134 706522
rect 364514 706202 364546 706438
rect 364782 706202 364866 706438
rect 365102 706202 365134 706438
rect 364514 691174 365134 706202
rect 364514 690938 364546 691174
rect 364782 690938 364866 691174
rect 365102 690938 365134 691174
rect 364514 690854 365134 690938
rect 364514 690618 364546 690854
rect 364782 690618 364866 690854
rect 365102 690618 365134 690854
rect 364514 655174 365134 690618
rect 364514 654938 364546 655174
rect 364782 654938 364866 655174
rect 365102 654938 365134 655174
rect 364514 654854 365134 654938
rect 364514 654618 364546 654854
rect 364782 654618 364866 654854
rect 365102 654618 365134 654854
rect 364514 619174 365134 654618
rect 364514 618938 364546 619174
rect 364782 618938 364866 619174
rect 365102 618938 365134 619174
rect 364514 618854 365134 618938
rect 364514 618618 364546 618854
rect 364782 618618 364866 618854
rect 365102 618618 365134 618854
rect 364514 583174 365134 618618
rect 364514 582938 364546 583174
rect 364782 582938 364866 583174
rect 365102 582938 365134 583174
rect 364514 582854 365134 582938
rect 364514 582618 364546 582854
rect 364782 582618 364866 582854
rect 365102 582618 365134 582854
rect 364514 547174 365134 582618
rect 364514 546938 364546 547174
rect 364782 546938 364866 547174
rect 365102 546938 365134 547174
rect 364514 546854 365134 546938
rect 364514 546618 364546 546854
rect 364782 546618 364866 546854
rect 365102 546618 365134 546854
rect 364514 511174 365134 546618
rect 364514 510938 364546 511174
rect 364782 510938 364866 511174
rect 365102 510938 365134 511174
rect 364514 510854 365134 510938
rect 364514 510618 364546 510854
rect 364782 510618 364866 510854
rect 365102 510618 365134 510854
rect 364514 475174 365134 510618
rect 364514 474938 364546 475174
rect 364782 474938 364866 475174
rect 365102 474938 365134 475174
rect 364514 474854 365134 474938
rect 364514 474618 364546 474854
rect 364782 474618 364866 474854
rect 365102 474618 365134 474854
rect 364514 439174 365134 474618
rect 364514 438938 364546 439174
rect 364782 438938 364866 439174
rect 365102 438938 365134 439174
rect 364514 438854 365134 438938
rect 364514 438618 364546 438854
rect 364782 438618 364866 438854
rect 365102 438618 365134 438854
rect 364514 403174 365134 438618
rect 364514 402938 364546 403174
rect 364782 402938 364866 403174
rect 365102 402938 365134 403174
rect 364514 402854 365134 402938
rect 364514 402618 364546 402854
rect 364782 402618 364866 402854
rect 365102 402618 365134 402854
rect 364514 367174 365134 402618
rect 364514 366938 364546 367174
rect 364782 366938 364866 367174
rect 365102 366938 365134 367174
rect 364514 366854 365134 366938
rect 364514 366618 364546 366854
rect 364782 366618 364866 366854
rect 365102 366618 365134 366854
rect 364514 331174 365134 366618
rect 364514 330938 364546 331174
rect 364782 330938 364866 331174
rect 365102 330938 365134 331174
rect 364514 330854 365134 330938
rect 364514 330618 364546 330854
rect 364782 330618 364866 330854
rect 365102 330618 365134 330854
rect 364514 295174 365134 330618
rect 364514 294938 364546 295174
rect 364782 294938 364866 295174
rect 365102 294938 365134 295174
rect 364514 294854 365134 294938
rect 364514 294618 364546 294854
rect 364782 294618 364866 294854
rect 365102 294618 365134 294854
rect 364514 259174 365134 294618
rect 364514 258938 364546 259174
rect 364782 258938 364866 259174
rect 365102 258938 365134 259174
rect 364514 258854 365134 258938
rect 364514 258618 364546 258854
rect 364782 258618 364866 258854
rect 365102 258618 365134 258854
rect 364514 223174 365134 258618
rect 364514 222938 364546 223174
rect 364782 222938 364866 223174
rect 365102 222938 365134 223174
rect 364514 222854 365134 222938
rect 364514 222618 364546 222854
rect 364782 222618 364866 222854
rect 365102 222618 365134 222854
rect 364514 187174 365134 222618
rect 364514 186938 364546 187174
rect 364782 186938 364866 187174
rect 365102 186938 365134 187174
rect 364514 186854 365134 186938
rect 364514 186618 364546 186854
rect 364782 186618 364866 186854
rect 365102 186618 365134 186854
rect 364514 151174 365134 186618
rect 364514 150938 364546 151174
rect 364782 150938 364866 151174
rect 365102 150938 365134 151174
rect 364514 150854 365134 150938
rect 364514 150618 364546 150854
rect 364782 150618 364866 150854
rect 365102 150618 365134 150854
rect 364514 115174 365134 150618
rect 364514 114938 364546 115174
rect 364782 114938 364866 115174
rect 365102 114938 365134 115174
rect 364514 114854 365134 114938
rect 364514 114618 364546 114854
rect 364782 114618 364866 114854
rect 365102 114618 365134 114854
rect 364514 79174 365134 114618
rect 364514 78938 364546 79174
rect 364782 78938 364866 79174
rect 365102 78938 365134 79174
rect 364514 78854 365134 78938
rect 364514 78618 364546 78854
rect 364782 78618 364866 78854
rect 365102 78618 365134 78854
rect 364514 43174 365134 78618
rect 364514 42938 364546 43174
rect 364782 42938 364866 43174
rect 365102 42938 365134 43174
rect 364514 42854 365134 42938
rect 364514 42618 364546 42854
rect 364782 42618 364866 42854
rect 365102 42618 365134 42854
rect 364514 7174 365134 42618
rect 364514 6938 364546 7174
rect 364782 6938 364866 7174
rect 365102 6938 365134 7174
rect 364514 6854 365134 6938
rect 364514 6618 364546 6854
rect 364782 6618 364866 6854
rect 365102 6618 365134 6854
rect 364514 -2266 365134 6618
rect 364514 -2502 364546 -2266
rect 364782 -2502 364866 -2266
rect 365102 -2502 365134 -2266
rect 364514 -2586 365134 -2502
rect 364514 -2822 364546 -2586
rect 364782 -2822 364866 -2586
rect 365102 -2822 365134 -2586
rect 364514 -3814 365134 -2822
rect 368234 694894 368854 708122
rect 368234 694658 368266 694894
rect 368502 694658 368586 694894
rect 368822 694658 368854 694894
rect 368234 694574 368854 694658
rect 368234 694338 368266 694574
rect 368502 694338 368586 694574
rect 368822 694338 368854 694574
rect 368234 658894 368854 694338
rect 368234 658658 368266 658894
rect 368502 658658 368586 658894
rect 368822 658658 368854 658894
rect 368234 658574 368854 658658
rect 368234 658338 368266 658574
rect 368502 658338 368586 658574
rect 368822 658338 368854 658574
rect 368234 622894 368854 658338
rect 368234 622658 368266 622894
rect 368502 622658 368586 622894
rect 368822 622658 368854 622894
rect 368234 622574 368854 622658
rect 368234 622338 368266 622574
rect 368502 622338 368586 622574
rect 368822 622338 368854 622574
rect 368234 586894 368854 622338
rect 368234 586658 368266 586894
rect 368502 586658 368586 586894
rect 368822 586658 368854 586894
rect 368234 586574 368854 586658
rect 368234 586338 368266 586574
rect 368502 586338 368586 586574
rect 368822 586338 368854 586574
rect 368234 550894 368854 586338
rect 368234 550658 368266 550894
rect 368502 550658 368586 550894
rect 368822 550658 368854 550894
rect 368234 550574 368854 550658
rect 368234 550338 368266 550574
rect 368502 550338 368586 550574
rect 368822 550338 368854 550574
rect 368234 514894 368854 550338
rect 368234 514658 368266 514894
rect 368502 514658 368586 514894
rect 368822 514658 368854 514894
rect 368234 514574 368854 514658
rect 368234 514338 368266 514574
rect 368502 514338 368586 514574
rect 368822 514338 368854 514574
rect 368234 478894 368854 514338
rect 368234 478658 368266 478894
rect 368502 478658 368586 478894
rect 368822 478658 368854 478894
rect 368234 478574 368854 478658
rect 368234 478338 368266 478574
rect 368502 478338 368586 478574
rect 368822 478338 368854 478574
rect 368234 442894 368854 478338
rect 368234 442658 368266 442894
rect 368502 442658 368586 442894
rect 368822 442658 368854 442894
rect 368234 442574 368854 442658
rect 368234 442338 368266 442574
rect 368502 442338 368586 442574
rect 368822 442338 368854 442574
rect 368234 406894 368854 442338
rect 368234 406658 368266 406894
rect 368502 406658 368586 406894
rect 368822 406658 368854 406894
rect 368234 406574 368854 406658
rect 368234 406338 368266 406574
rect 368502 406338 368586 406574
rect 368822 406338 368854 406574
rect 368234 370894 368854 406338
rect 368234 370658 368266 370894
rect 368502 370658 368586 370894
rect 368822 370658 368854 370894
rect 368234 370574 368854 370658
rect 368234 370338 368266 370574
rect 368502 370338 368586 370574
rect 368822 370338 368854 370574
rect 368234 334894 368854 370338
rect 368234 334658 368266 334894
rect 368502 334658 368586 334894
rect 368822 334658 368854 334894
rect 368234 334574 368854 334658
rect 368234 334338 368266 334574
rect 368502 334338 368586 334574
rect 368822 334338 368854 334574
rect 368234 298894 368854 334338
rect 368234 298658 368266 298894
rect 368502 298658 368586 298894
rect 368822 298658 368854 298894
rect 368234 298574 368854 298658
rect 368234 298338 368266 298574
rect 368502 298338 368586 298574
rect 368822 298338 368854 298574
rect 368234 262894 368854 298338
rect 368234 262658 368266 262894
rect 368502 262658 368586 262894
rect 368822 262658 368854 262894
rect 368234 262574 368854 262658
rect 368234 262338 368266 262574
rect 368502 262338 368586 262574
rect 368822 262338 368854 262574
rect 368234 226894 368854 262338
rect 368234 226658 368266 226894
rect 368502 226658 368586 226894
rect 368822 226658 368854 226894
rect 368234 226574 368854 226658
rect 368234 226338 368266 226574
rect 368502 226338 368586 226574
rect 368822 226338 368854 226574
rect 368234 190894 368854 226338
rect 368234 190658 368266 190894
rect 368502 190658 368586 190894
rect 368822 190658 368854 190894
rect 368234 190574 368854 190658
rect 368234 190338 368266 190574
rect 368502 190338 368586 190574
rect 368822 190338 368854 190574
rect 368234 154894 368854 190338
rect 368234 154658 368266 154894
rect 368502 154658 368586 154894
rect 368822 154658 368854 154894
rect 368234 154574 368854 154658
rect 368234 154338 368266 154574
rect 368502 154338 368586 154574
rect 368822 154338 368854 154574
rect 368234 118894 368854 154338
rect 368234 118658 368266 118894
rect 368502 118658 368586 118894
rect 368822 118658 368854 118894
rect 368234 118574 368854 118658
rect 368234 118338 368266 118574
rect 368502 118338 368586 118574
rect 368822 118338 368854 118574
rect 368234 82894 368854 118338
rect 368234 82658 368266 82894
rect 368502 82658 368586 82894
rect 368822 82658 368854 82894
rect 368234 82574 368854 82658
rect 368234 82338 368266 82574
rect 368502 82338 368586 82574
rect 368822 82338 368854 82574
rect 368234 46894 368854 82338
rect 368234 46658 368266 46894
rect 368502 46658 368586 46894
rect 368822 46658 368854 46894
rect 368234 46574 368854 46658
rect 368234 46338 368266 46574
rect 368502 46338 368586 46574
rect 368822 46338 368854 46574
rect 368234 10894 368854 46338
rect 368234 10658 368266 10894
rect 368502 10658 368586 10894
rect 368822 10658 368854 10894
rect 368234 10574 368854 10658
rect 368234 10338 368266 10574
rect 368502 10338 368586 10574
rect 368822 10338 368854 10574
rect 368234 -4186 368854 10338
rect 370794 705798 371414 705830
rect 370794 705562 370826 705798
rect 371062 705562 371146 705798
rect 371382 705562 371414 705798
rect 370794 705478 371414 705562
rect 370794 705242 370826 705478
rect 371062 705242 371146 705478
rect 371382 705242 371414 705478
rect 370794 669454 371414 705242
rect 370794 669218 370826 669454
rect 371062 669218 371146 669454
rect 371382 669218 371414 669454
rect 370794 669134 371414 669218
rect 370794 668898 370826 669134
rect 371062 668898 371146 669134
rect 371382 668898 371414 669134
rect 370794 633454 371414 668898
rect 370794 633218 370826 633454
rect 371062 633218 371146 633454
rect 371382 633218 371414 633454
rect 370794 633134 371414 633218
rect 370794 632898 370826 633134
rect 371062 632898 371146 633134
rect 371382 632898 371414 633134
rect 370794 597454 371414 632898
rect 370794 597218 370826 597454
rect 371062 597218 371146 597454
rect 371382 597218 371414 597454
rect 370794 597134 371414 597218
rect 370794 596898 370826 597134
rect 371062 596898 371146 597134
rect 371382 596898 371414 597134
rect 370794 561454 371414 596898
rect 370794 561218 370826 561454
rect 371062 561218 371146 561454
rect 371382 561218 371414 561454
rect 370794 561134 371414 561218
rect 370794 560898 370826 561134
rect 371062 560898 371146 561134
rect 371382 560898 371414 561134
rect 370794 525454 371414 560898
rect 370794 525218 370826 525454
rect 371062 525218 371146 525454
rect 371382 525218 371414 525454
rect 370794 525134 371414 525218
rect 370794 524898 370826 525134
rect 371062 524898 371146 525134
rect 371382 524898 371414 525134
rect 370794 489454 371414 524898
rect 370794 489218 370826 489454
rect 371062 489218 371146 489454
rect 371382 489218 371414 489454
rect 370794 489134 371414 489218
rect 370794 488898 370826 489134
rect 371062 488898 371146 489134
rect 371382 488898 371414 489134
rect 370794 453454 371414 488898
rect 370794 453218 370826 453454
rect 371062 453218 371146 453454
rect 371382 453218 371414 453454
rect 370794 453134 371414 453218
rect 370794 452898 370826 453134
rect 371062 452898 371146 453134
rect 371382 452898 371414 453134
rect 370794 417454 371414 452898
rect 370794 417218 370826 417454
rect 371062 417218 371146 417454
rect 371382 417218 371414 417454
rect 370794 417134 371414 417218
rect 370794 416898 370826 417134
rect 371062 416898 371146 417134
rect 371382 416898 371414 417134
rect 370794 381454 371414 416898
rect 370794 381218 370826 381454
rect 371062 381218 371146 381454
rect 371382 381218 371414 381454
rect 370794 381134 371414 381218
rect 370794 380898 370826 381134
rect 371062 380898 371146 381134
rect 371382 380898 371414 381134
rect 370794 345454 371414 380898
rect 370794 345218 370826 345454
rect 371062 345218 371146 345454
rect 371382 345218 371414 345454
rect 370794 345134 371414 345218
rect 370794 344898 370826 345134
rect 371062 344898 371146 345134
rect 371382 344898 371414 345134
rect 370794 309454 371414 344898
rect 370794 309218 370826 309454
rect 371062 309218 371146 309454
rect 371382 309218 371414 309454
rect 370794 309134 371414 309218
rect 370794 308898 370826 309134
rect 371062 308898 371146 309134
rect 371382 308898 371414 309134
rect 370794 273454 371414 308898
rect 370794 273218 370826 273454
rect 371062 273218 371146 273454
rect 371382 273218 371414 273454
rect 370794 273134 371414 273218
rect 370794 272898 370826 273134
rect 371062 272898 371146 273134
rect 371382 272898 371414 273134
rect 370794 237454 371414 272898
rect 370794 237218 370826 237454
rect 371062 237218 371146 237454
rect 371382 237218 371414 237454
rect 370794 237134 371414 237218
rect 370794 236898 370826 237134
rect 371062 236898 371146 237134
rect 371382 236898 371414 237134
rect 370794 201454 371414 236898
rect 370794 201218 370826 201454
rect 371062 201218 371146 201454
rect 371382 201218 371414 201454
rect 370794 201134 371414 201218
rect 370794 200898 370826 201134
rect 371062 200898 371146 201134
rect 371382 200898 371414 201134
rect 370794 165454 371414 200898
rect 370794 165218 370826 165454
rect 371062 165218 371146 165454
rect 371382 165218 371414 165454
rect 370794 165134 371414 165218
rect 370794 164898 370826 165134
rect 371062 164898 371146 165134
rect 371382 164898 371414 165134
rect 370794 129454 371414 164898
rect 370794 129218 370826 129454
rect 371062 129218 371146 129454
rect 371382 129218 371414 129454
rect 370794 129134 371414 129218
rect 370794 128898 370826 129134
rect 371062 128898 371146 129134
rect 371382 128898 371414 129134
rect 370794 93454 371414 128898
rect 370794 93218 370826 93454
rect 371062 93218 371146 93454
rect 371382 93218 371414 93454
rect 370794 93134 371414 93218
rect 370794 92898 370826 93134
rect 371062 92898 371146 93134
rect 371382 92898 371414 93134
rect 370794 57454 371414 92898
rect 370794 57218 370826 57454
rect 371062 57218 371146 57454
rect 371382 57218 371414 57454
rect 370794 57134 371414 57218
rect 370794 56898 370826 57134
rect 371062 56898 371146 57134
rect 371382 56898 371414 57134
rect 370794 21454 371414 56898
rect 370794 21218 370826 21454
rect 371062 21218 371146 21454
rect 371382 21218 371414 21454
rect 370794 21134 371414 21218
rect 370794 20898 370826 21134
rect 371062 20898 371146 21134
rect 371382 20898 371414 21134
rect 370794 -1306 371414 20898
rect 370794 -1542 370826 -1306
rect 371062 -1542 371146 -1306
rect 371382 -1542 371414 -1306
rect 370794 -1626 371414 -1542
rect 370794 -1862 370826 -1626
rect 371062 -1862 371146 -1626
rect 371382 -1862 371414 -1626
rect 370794 -1894 371414 -1862
rect 371954 698614 372574 710042
rect 381954 711558 382574 711590
rect 381954 711322 381986 711558
rect 382222 711322 382306 711558
rect 382542 711322 382574 711558
rect 381954 711238 382574 711322
rect 381954 711002 381986 711238
rect 382222 711002 382306 711238
rect 382542 711002 382574 711238
rect 378234 709638 378854 709670
rect 378234 709402 378266 709638
rect 378502 709402 378586 709638
rect 378822 709402 378854 709638
rect 378234 709318 378854 709402
rect 378234 709082 378266 709318
rect 378502 709082 378586 709318
rect 378822 709082 378854 709318
rect 371954 698378 371986 698614
rect 372222 698378 372306 698614
rect 372542 698378 372574 698614
rect 371954 698294 372574 698378
rect 371954 698058 371986 698294
rect 372222 698058 372306 698294
rect 372542 698058 372574 698294
rect 371954 662614 372574 698058
rect 371954 662378 371986 662614
rect 372222 662378 372306 662614
rect 372542 662378 372574 662614
rect 371954 662294 372574 662378
rect 371954 662058 371986 662294
rect 372222 662058 372306 662294
rect 372542 662058 372574 662294
rect 371954 626614 372574 662058
rect 371954 626378 371986 626614
rect 372222 626378 372306 626614
rect 372542 626378 372574 626614
rect 371954 626294 372574 626378
rect 371954 626058 371986 626294
rect 372222 626058 372306 626294
rect 372542 626058 372574 626294
rect 371954 590614 372574 626058
rect 371954 590378 371986 590614
rect 372222 590378 372306 590614
rect 372542 590378 372574 590614
rect 371954 590294 372574 590378
rect 371954 590058 371986 590294
rect 372222 590058 372306 590294
rect 372542 590058 372574 590294
rect 371954 554614 372574 590058
rect 371954 554378 371986 554614
rect 372222 554378 372306 554614
rect 372542 554378 372574 554614
rect 371954 554294 372574 554378
rect 371954 554058 371986 554294
rect 372222 554058 372306 554294
rect 372542 554058 372574 554294
rect 371954 518614 372574 554058
rect 371954 518378 371986 518614
rect 372222 518378 372306 518614
rect 372542 518378 372574 518614
rect 371954 518294 372574 518378
rect 371954 518058 371986 518294
rect 372222 518058 372306 518294
rect 372542 518058 372574 518294
rect 371954 482614 372574 518058
rect 371954 482378 371986 482614
rect 372222 482378 372306 482614
rect 372542 482378 372574 482614
rect 371954 482294 372574 482378
rect 371954 482058 371986 482294
rect 372222 482058 372306 482294
rect 372542 482058 372574 482294
rect 371954 446614 372574 482058
rect 371954 446378 371986 446614
rect 372222 446378 372306 446614
rect 372542 446378 372574 446614
rect 371954 446294 372574 446378
rect 371954 446058 371986 446294
rect 372222 446058 372306 446294
rect 372542 446058 372574 446294
rect 371954 410614 372574 446058
rect 371954 410378 371986 410614
rect 372222 410378 372306 410614
rect 372542 410378 372574 410614
rect 371954 410294 372574 410378
rect 371954 410058 371986 410294
rect 372222 410058 372306 410294
rect 372542 410058 372574 410294
rect 371954 374614 372574 410058
rect 371954 374378 371986 374614
rect 372222 374378 372306 374614
rect 372542 374378 372574 374614
rect 371954 374294 372574 374378
rect 371954 374058 371986 374294
rect 372222 374058 372306 374294
rect 372542 374058 372574 374294
rect 371954 338614 372574 374058
rect 371954 338378 371986 338614
rect 372222 338378 372306 338614
rect 372542 338378 372574 338614
rect 371954 338294 372574 338378
rect 371954 338058 371986 338294
rect 372222 338058 372306 338294
rect 372542 338058 372574 338294
rect 371954 302614 372574 338058
rect 371954 302378 371986 302614
rect 372222 302378 372306 302614
rect 372542 302378 372574 302614
rect 371954 302294 372574 302378
rect 371954 302058 371986 302294
rect 372222 302058 372306 302294
rect 372542 302058 372574 302294
rect 371954 266614 372574 302058
rect 371954 266378 371986 266614
rect 372222 266378 372306 266614
rect 372542 266378 372574 266614
rect 371954 266294 372574 266378
rect 371954 266058 371986 266294
rect 372222 266058 372306 266294
rect 372542 266058 372574 266294
rect 371954 230614 372574 266058
rect 371954 230378 371986 230614
rect 372222 230378 372306 230614
rect 372542 230378 372574 230614
rect 371954 230294 372574 230378
rect 371954 230058 371986 230294
rect 372222 230058 372306 230294
rect 372542 230058 372574 230294
rect 371954 194614 372574 230058
rect 371954 194378 371986 194614
rect 372222 194378 372306 194614
rect 372542 194378 372574 194614
rect 371954 194294 372574 194378
rect 371954 194058 371986 194294
rect 372222 194058 372306 194294
rect 372542 194058 372574 194294
rect 371954 158614 372574 194058
rect 371954 158378 371986 158614
rect 372222 158378 372306 158614
rect 372542 158378 372574 158614
rect 371954 158294 372574 158378
rect 371954 158058 371986 158294
rect 372222 158058 372306 158294
rect 372542 158058 372574 158294
rect 371954 122614 372574 158058
rect 371954 122378 371986 122614
rect 372222 122378 372306 122614
rect 372542 122378 372574 122614
rect 371954 122294 372574 122378
rect 371954 122058 371986 122294
rect 372222 122058 372306 122294
rect 372542 122058 372574 122294
rect 371954 86614 372574 122058
rect 371954 86378 371986 86614
rect 372222 86378 372306 86614
rect 372542 86378 372574 86614
rect 371954 86294 372574 86378
rect 371954 86058 371986 86294
rect 372222 86058 372306 86294
rect 372542 86058 372574 86294
rect 371954 50614 372574 86058
rect 371954 50378 371986 50614
rect 372222 50378 372306 50614
rect 372542 50378 372574 50614
rect 371954 50294 372574 50378
rect 371954 50058 371986 50294
rect 372222 50058 372306 50294
rect 372542 50058 372574 50294
rect 371954 14614 372574 50058
rect 371954 14378 371986 14614
rect 372222 14378 372306 14614
rect 372542 14378 372574 14614
rect 371954 14294 372574 14378
rect 371954 14058 371986 14294
rect 372222 14058 372306 14294
rect 372542 14058 372574 14294
rect 368234 -4422 368266 -4186
rect 368502 -4422 368586 -4186
rect 368822 -4422 368854 -4186
rect 368234 -4506 368854 -4422
rect 368234 -4742 368266 -4506
rect 368502 -4742 368586 -4506
rect 368822 -4742 368854 -4506
rect 368234 -5734 368854 -4742
rect 361954 -7302 361986 -7066
rect 362222 -7302 362306 -7066
rect 362542 -7302 362574 -7066
rect 361954 -7386 362574 -7302
rect 361954 -7622 361986 -7386
rect 362222 -7622 362306 -7386
rect 362542 -7622 362574 -7386
rect 361954 -7654 362574 -7622
rect 371954 -6106 372574 14058
rect 374514 707718 375134 707750
rect 374514 707482 374546 707718
rect 374782 707482 374866 707718
rect 375102 707482 375134 707718
rect 374514 707398 375134 707482
rect 374514 707162 374546 707398
rect 374782 707162 374866 707398
rect 375102 707162 375134 707398
rect 374514 673174 375134 707162
rect 374514 672938 374546 673174
rect 374782 672938 374866 673174
rect 375102 672938 375134 673174
rect 374514 672854 375134 672938
rect 374514 672618 374546 672854
rect 374782 672618 374866 672854
rect 375102 672618 375134 672854
rect 374514 637174 375134 672618
rect 374514 636938 374546 637174
rect 374782 636938 374866 637174
rect 375102 636938 375134 637174
rect 374514 636854 375134 636938
rect 374514 636618 374546 636854
rect 374782 636618 374866 636854
rect 375102 636618 375134 636854
rect 374514 601174 375134 636618
rect 374514 600938 374546 601174
rect 374782 600938 374866 601174
rect 375102 600938 375134 601174
rect 374514 600854 375134 600938
rect 374514 600618 374546 600854
rect 374782 600618 374866 600854
rect 375102 600618 375134 600854
rect 374514 565174 375134 600618
rect 374514 564938 374546 565174
rect 374782 564938 374866 565174
rect 375102 564938 375134 565174
rect 374514 564854 375134 564938
rect 374514 564618 374546 564854
rect 374782 564618 374866 564854
rect 375102 564618 375134 564854
rect 374514 529174 375134 564618
rect 374514 528938 374546 529174
rect 374782 528938 374866 529174
rect 375102 528938 375134 529174
rect 374514 528854 375134 528938
rect 374514 528618 374546 528854
rect 374782 528618 374866 528854
rect 375102 528618 375134 528854
rect 374514 493174 375134 528618
rect 374514 492938 374546 493174
rect 374782 492938 374866 493174
rect 375102 492938 375134 493174
rect 374514 492854 375134 492938
rect 374514 492618 374546 492854
rect 374782 492618 374866 492854
rect 375102 492618 375134 492854
rect 374514 457174 375134 492618
rect 374514 456938 374546 457174
rect 374782 456938 374866 457174
rect 375102 456938 375134 457174
rect 374514 456854 375134 456938
rect 374514 456618 374546 456854
rect 374782 456618 374866 456854
rect 375102 456618 375134 456854
rect 374514 421174 375134 456618
rect 374514 420938 374546 421174
rect 374782 420938 374866 421174
rect 375102 420938 375134 421174
rect 374514 420854 375134 420938
rect 374514 420618 374546 420854
rect 374782 420618 374866 420854
rect 375102 420618 375134 420854
rect 374514 385174 375134 420618
rect 374514 384938 374546 385174
rect 374782 384938 374866 385174
rect 375102 384938 375134 385174
rect 374514 384854 375134 384938
rect 374514 384618 374546 384854
rect 374782 384618 374866 384854
rect 375102 384618 375134 384854
rect 374514 349174 375134 384618
rect 374514 348938 374546 349174
rect 374782 348938 374866 349174
rect 375102 348938 375134 349174
rect 374514 348854 375134 348938
rect 374514 348618 374546 348854
rect 374782 348618 374866 348854
rect 375102 348618 375134 348854
rect 374514 313174 375134 348618
rect 374514 312938 374546 313174
rect 374782 312938 374866 313174
rect 375102 312938 375134 313174
rect 374514 312854 375134 312938
rect 374514 312618 374546 312854
rect 374782 312618 374866 312854
rect 375102 312618 375134 312854
rect 374514 277174 375134 312618
rect 374514 276938 374546 277174
rect 374782 276938 374866 277174
rect 375102 276938 375134 277174
rect 374514 276854 375134 276938
rect 374514 276618 374546 276854
rect 374782 276618 374866 276854
rect 375102 276618 375134 276854
rect 374514 241174 375134 276618
rect 374514 240938 374546 241174
rect 374782 240938 374866 241174
rect 375102 240938 375134 241174
rect 374514 240854 375134 240938
rect 374514 240618 374546 240854
rect 374782 240618 374866 240854
rect 375102 240618 375134 240854
rect 374514 205174 375134 240618
rect 374514 204938 374546 205174
rect 374782 204938 374866 205174
rect 375102 204938 375134 205174
rect 374514 204854 375134 204938
rect 374514 204618 374546 204854
rect 374782 204618 374866 204854
rect 375102 204618 375134 204854
rect 374514 169174 375134 204618
rect 374514 168938 374546 169174
rect 374782 168938 374866 169174
rect 375102 168938 375134 169174
rect 374514 168854 375134 168938
rect 374514 168618 374546 168854
rect 374782 168618 374866 168854
rect 375102 168618 375134 168854
rect 374514 133174 375134 168618
rect 374514 132938 374546 133174
rect 374782 132938 374866 133174
rect 375102 132938 375134 133174
rect 374514 132854 375134 132938
rect 374514 132618 374546 132854
rect 374782 132618 374866 132854
rect 375102 132618 375134 132854
rect 374514 97174 375134 132618
rect 374514 96938 374546 97174
rect 374782 96938 374866 97174
rect 375102 96938 375134 97174
rect 374514 96854 375134 96938
rect 374514 96618 374546 96854
rect 374782 96618 374866 96854
rect 375102 96618 375134 96854
rect 374514 61174 375134 96618
rect 374514 60938 374546 61174
rect 374782 60938 374866 61174
rect 375102 60938 375134 61174
rect 374514 60854 375134 60938
rect 374514 60618 374546 60854
rect 374782 60618 374866 60854
rect 375102 60618 375134 60854
rect 374514 25174 375134 60618
rect 374514 24938 374546 25174
rect 374782 24938 374866 25174
rect 375102 24938 375134 25174
rect 374514 24854 375134 24938
rect 374514 24618 374546 24854
rect 374782 24618 374866 24854
rect 375102 24618 375134 24854
rect 374514 -3226 375134 24618
rect 374514 -3462 374546 -3226
rect 374782 -3462 374866 -3226
rect 375102 -3462 375134 -3226
rect 374514 -3546 375134 -3462
rect 374514 -3782 374546 -3546
rect 374782 -3782 374866 -3546
rect 375102 -3782 375134 -3546
rect 374514 -3814 375134 -3782
rect 378234 676894 378854 709082
rect 378234 676658 378266 676894
rect 378502 676658 378586 676894
rect 378822 676658 378854 676894
rect 378234 676574 378854 676658
rect 378234 676338 378266 676574
rect 378502 676338 378586 676574
rect 378822 676338 378854 676574
rect 378234 640894 378854 676338
rect 378234 640658 378266 640894
rect 378502 640658 378586 640894
rect 378822 640658 378854 640894
rect 378234 640574 378854 640658
rect 378234 640338 378266 640574
rect 378502 640338 378586 640574
rect 378822 640338 378854 640574
rect 378234 604894 378854 640338
rect 378234 604658 378266 604894
rect 378502 604658 378586 604894
rect 378822 604658 378854 604894
rect 378234 604574 378854 604658
rect 378234 604338 378266 604574
rect 378502 604338 378586 604574
rect 378822 604338 378854 604574
rect 378234 568894 378854 604338
rect 378234 568658 378266 568894
rect 378502 568658 378586 568894
rect 378822 568658 378854 568894
rect 378234 568574 378854 568658
rect 378234 568338 378266 568574
rect 378502 568338 378586 568574
rect 378822 568338 378854 568574
rect 378234 532894 378854 568338
rect 378234 532658 378266 532894
rect 378502 532658 378586 532894
rect 378822 532658 378854 532894
rect 378234 532574 378854 532658
rect 378234 532338 378266 532574
rect 378502 532338 378586 532574
rect 378822 532338 378854 532574
rect 378234 496894 378854 532338
rect 378234 496658 378266 496894
rect 378502 496658 378586 496894
rect 378822 496658 378854 496894
rect 378234 496574 378854 496658
rect 378234 496338 378266 496574
rect 378502 496338 378586 496574
rect 378822 496338 378854 496574
rect 378234 460894 378854 496338
rect 378234 460658 378266 460894
rect 378502 460658 378586 460894
rect 378822 460658 378854 460894
rect 378234 460574 378854 460658
rect 378234 460338 378266 460574
rect 378502 460338 378586 460574
rect 378822 460338 378854 460574
rect 378234 424894 378854 460338
rect 378234 424658 378266 424894
rect 378502 424658 378586 424894
rect 378822 424658 378854 424894
rect 378234 424574 378854 424658
rect 378234 424338 378266 424574
rect 378502 424338 378586 424574
rect 378822 424338 378854 424574
rect 378234 388894 378854 424338
rect 378234 388658 378266 388894
rect 378502 388658 378586 388894
rect 378822 388658 378854 388894
rect 378234 388574 378854 388658
rect 378234 388338 378266 388574
rect 378502 388338 378586 388574
rect 378822 388338 378854 388574
rect 378234 352894 378854 388338
rect 378234 352658 378266 352894
rect 378502 352658 378586 352894
rect 378822 352658 378854 352894
rect 378234 352574 378854 352658
rect 378234 352338 378266 352574
rect 378502 352338 378586 352574
rect 378822 352338 378854 352574
rect 378234 316894 378854 352338
rect 378234 316658 378266 316894
rect 378502 316658 378586 316894
rect 378822 316658 378854 316894
rect 378234 316574 378854 316658
rect 378234 316338 378266 316574
rect 378502 316338 378586 316574
rect 378822 316338 378854 316574
rect 378234 280894 378854 316338
rect 378234 280658 378266 280894
rect 378502 280658 378586 280894
rect 378822 280658 378854 280894
rect 378234 280574 378854 280658
rect 378234 280338 378266 280574
rect 378502 280338 378586 280574
rect 378822 280338 378854 280574
rect 378234 244894 378854 280338
rect 378234 244658 378266 244894
rect 378502 244658 378586 244894
rect 378822 244658 378854 244894
rect 378234 244574 378854 244658
rect 378234 244338 378266 244574
rect 378502 244338 378586 244574
rect 378822 244338 378854 244574
rect 378234 208894 378854 244338
rect 378234 208658 378266 208894
rect 378502 208658 378586 208894
rect 378822 208658 378854 208894
rect 378234 208574 378854 208658
rect 378234 208338 378266 208574
rect 378502 208338 378586 208574
rect 378822 208338 378854 208574
rect 378234 172894 378854 208338
rect 378234 172658 378266 172894
rect 378502 172658 378586 172894
rect 378822 172658 378854 172894
rect 378234 172574 378854 172658
rect 378234 172338 378266 172574
rect 378502 172338 378586 172574
rect 378822 172338 378854 172574
rect 378234 136894 378854 172338
rect 378234 136658 378266 136894
rect 378502 136658 378586 136894
rect 378822 136658 378854 136894
rect 378234 136574 378854 136658
rect 378234 136338 378266 136574
rect 378502 136338 378586 136574
rect 378822 136338 378854 136574
rect 378234 100894 378854 136338
rect 378234 100658 378266 100894
rect 378502 100658 378586 100894
rect 378822 100658 378854 100894
rect 378234 100574 378854 100658
rect 378234 100338 378266 100574
rect 378502 100338 378586 100574
rect 378822 100338 378854 100574
rect 378234 64894 378854 100338
rect 378234 64658 378266 64894
rect 378502 64658 378586 64894
rect 378822 64658 378854 64894
rect 378234 64574 378854 64658
rect 378234 64338 378266 64574
rect 378502 64338 378586 64574
rect 378822 64338 378854 64574
rect 378234 28894 378854 64338
rect 378234 28658 378266 28894
rect 378502 28658 378586 28894
rect 378822 28658 378854 28894
rect 378234 28574 378854 28658
rect 378234 28338 378266 28574
rect 378502 28338 378586 28574
rect 378822 28338 378854 28574
rect 378234 -5146 378854 28338
rect 380794 704838 381414 705830
rect 380794 704602 380826 704838
rect 381062 704602 381146 704838
rect 381382 704602 381414 704838
rect 380794 704518 381414 704602
rect 380794 704282 380826 704518
rect 381062 704282 381146 704518
rect 381382 704282 381414 704518
rect 380794 687454 381414 704282
rect 380794 687218 380826 687454
rect 381062 687218 381146 687454
rect 381382 687218 381414 687454
rect 380794 687134 381414 687218
rect 380794 686898 380826 687134
rect 381062 686898 381146 687134
rect 381382 686898 381414 687134
rect 380794 651454 381414 686898
rect 380794 651218 380826 651454
rect 381062 651218 381146 651454
rect 381382 651218 381414 651454
rect 380794 651134 381414 651218
rect 380794 650898 380826 651134
rect 381062 650898 381146 651134
rect 381382 650898 381414 651134
rect 380794 615454 381414 650898
rect 380794 615218 380826 615454
rect 381062 615218 381146 615454
rect 381382 615218 381414 615454
rect 380794 615134 381414 615218
rect 380794 614898 380826 615134
rect 381062 614898 381146 615134
rect 381382 614898 381414 615134
rect 380794 579454 381414 614898
rect 380794 579218 380826 579454
rect 381062 579218 381146 579454
rect 381382 579218 381414 579454
rect 380794 579134 381414 579218
rect 380794 578898 380826 579134
rect 381062 578898 381146 579134
rect 381382 578898 381414 579134
rect 380794 543454 381414 578898
rect 380794 543218 380826 543454
rect 381062 543218 381146 543454
rect 381382 543218 381414 543454
rect 380794 543134 381414 543218
rect 380794 542898 380826 543134
rect 381062 542898 381146 543134
rect 381382 542898 381414 543134
rect 380794 507454 381414 542898
rect 380794 507218 380826 507454
rect 381062 507218 381146 507454
rect 381382 507218 381414 507454
rect 380794 507134 381414 507218
rect 380794 506898 380826 507134
rect 381062 506898 381146 507134
rect 381382 506898 381414 507134
rect 380794 471454 381414 506898
rect 380794 471218 380826 471454
rect 381062 471218 381146 471454
rect 381382 471218 381414 471454
rect 380794 471134 381414 471218
rect 380794 470898 380826 471134
rect 381062 470898 381146 471134
rect 381382 470898 381414 471134
rect 380794 435454 381414 470898
rect 380794 435218 380826 435454
rect 381062 435218 381146 435454
rect 381382 435218 381414 435454
rect 380794 435134 381414 435218
rect 380794 434898 380826 435134
rect 381062 434898 381146 435134
rect 381382 434898 381414 435134
rect 380794 399454 381414 434898
rect 380794 399218 380826 399454
rect 381062 399218 381146 399454
rect 381382 399218 381414 399454
rect 380794 399134 381414 399218
rect 380794 398898 380826 399134
rect 381062 398898 381146 399134
rect 381382 398898 381414 399134
rect 380794 363454 381414 398898
rect 380794 363218 380826 363454
rect 381062 363218 381146 363454
rect 381382 363218 381414 363454
rect 380794 363134 381414 363218
rect 380794 362898 380826 363134
rect 381062 362898 381146 363134
rect 381382 362898 381414 363134
rect 380794 327454 381414 362898
rect 380794 327218 380826 327454
rect 381062 327218 381146 327454
rect 381382 327218 381414 327454
rect 380794 327134 381414 327218
rect 380794 326898 380826 327134
rect 381062 326898 381146 327134
rect 381382 326898 381414 327134
rect 380794 291454 381414 326898
rect 380794 291218 380826 291454
rect 381062 291218 381146 291454
rect 381382 291218 381414 291454
rect 380794 291134 381414 291218
rect 380794 290898 380826 291134
rect 381062 290898 381146 291134
rect 381382 290898 381414 291134
rect 380794 255454 381414 290898
rect 380794 255218 380826 255454
rect 381062 255218 381146 255454
rect 381382 255218 381414 255454
rect 380794 255134 381414 255218
rect 380794 254898 380826 255134
rect 381062 254898 381146 255134
rect 381382 254898 381414 255134
rect 380794 219454 381414 254898
rect 380794 219218 380826 219454
rect 381062 219218 381146 219454
rect 381382 219218 381414 219454
rect 380794 219134 381414 219218
rect 380794 218898 380826 219134
rect 381062 218898 381146 219134
rect 381382 218898 381414 219134
rect 380794 183454 381414 218898
rect 380794 183218 380826 183454
rect 381062 183218 381146 183454
rect 381382 183218 381414 183454
rect 380794 183134 381414 183218
rect 380794 182898 380826 183134
rect 381062 182898 381146 183134
rect 381382 182898 381414 183134
rect 380794 147454 381414 182898
rect 380794 147218 380826 147454
rect 381062 147218 381146 147454
rect 381382 147218 381414 147454
rect 380794 147134 381414 147218
rect 380794 146898 380826 147134
rect 381062 146898 381146 147134
rect 381382 146898 381414 147134
rect 380794 111454 381414 146898
rect 380794 111218 380826 111454
rect 381062 111218 381146 111454
rect 381382 111218 381414 111454
rect 380794 111134 381414 111218
rect 380794 110898 380826 111134
rect 381062 110898 381146 111134
rect 381382 110898 381414 111134
rect 380794 75454 381414 110898
rect 380794 75218 380826 75454
rect 381062 75218 381146 75454
rect 381382 75218 381414 75454
rect 380794 75134 381414 75218
rect 380794 74898 380826 75134
rect 381062 74898 381146 75134
rect 381382 74898 381414 75134
rect 380794 39454 381414 74898
rect 380794 39218 380826 39454
rect 381062 39218 381146 39454
rect 381382 39218 381414 39454
rect 380794 39134 381414 39218
rect 380794 38898 380826 39134
rect 381062 38898 381146 39134
rect 381382 38898 381414 39134
rect 380794 3454 381414 38898
rect 380794 3218 380826 3454
rect 381062 3218 381146 3454
rect 381382 3218 381414 3454
rect 380794 3134 381414 3218
rect 380794 2898 380826 3134
rect 381062 2898 381146 3134
rect 381382 2898 381414 3134
rect 380794 -346 381414 2898
rect 380794 -582 380826 -346
rect 381062 -582 381146 -346
rect 381382 -582 381414 -346
rect 380794 -666 381414 -582
rect 380794 -902 380826 -666
rect 381062 -902 381146 -666
rect 381382 -902 381414 -666
rect 380794 -1894 381414 -902
rect 381954 680614 382574 711002
rect 391954 710598 392574 711590
rect 391954 710362 391986 710598
rect 392222 710362 392306 710598
rect 392542 710362 392574 710598
rect 391954 710278 392574 710362
rect 391954 710042 391986 710278
rect 392222 710042 392306 710278
rect 392542 710042 392574 710278
rect 388234 708678 388854 709670
rect 388234 708442 388266 708678
rect 388502 708442 388586 708678
rect 388822 708442 388854 708678
rect 388234 708358 388854 708442
rect 388234 708122 388266 708358
rect 388502 708122 388586 708358
rect 388822 708122 388854 708358
rect 381954 680378 381986 680614
rect 382222 680378 382306 680614
rect 382542 680378 382574 680614
rect 381954 680294 382574 680378
rect 381954 680058 381986 680294
rect 382222 680058 382306 680294
rect 382542 680058 382574 680294
rect 381954 644614 382574 680058
rect 381954 644378 381986 644614
rect 382222 644378 382306 644614
rect 382542 644378 382574 644614
rect 381954 644294 382574 644378
rect 381954 644058 381986 644294
rect 382222 644058 382306 644294
rect 382542 644058 382574 644294
rect 381954 608614 382574 644058
rect 381954 608378 381986 608614
rect 382222 608378 382306 608614
rect 382542 608378 382574 608614
rect 381954 608294 382574 608378
rect 381954 608058 381986 608294
rect 382222 608058 382306 608294
rect 382542 608058 382574 608294
rect 381954 572614 382574 608058
rect 381954 572378 381986 572614
rect 382222 572378 382306 572614
rect 382542 572378 382574 572614
rect 381954 572294 382574 572378
rect 381954 572058 381986 572294
rect 382222 572058 382306 572294
rect 382542 572058 382574 572294
rect 381954 536614 382574 572058
rect 381954 536378 381986 536614
rect 382222 536378 382306 536614
rect 382542 536378 382574 536614
rect 381954 536294 382574 536378
rect 381954 536058 381986 536294
rect 382222 536058 382306 536294
rect 382542 536058 382574 536294
rect 381954 500614 382574 536058
rect 381954 500378 381986 500614
rect 382222 500378 382306 500614
rect 382542 500378 382574 500614
rect 381954 500294 382574 500378
rect 381954 500058 381986 500294
rect 382222 500058 382306 500294
rect 382542 500058 382574 500294
rect 381954 464614 382574 500058
rect 381954 464378 381986 464614
rect 382222 464378 382306 464614
rect 382542 464378 382574 464614
rect 381954 464294 382574 464378
rect 381954 464058 381986 464294
rect 382222 464058 382306 464294
rect 382542 464058 382574 464294
rect 381954 428614 382574 464058
rect 381954 428378 381986 428614
rect 382222 428378 382306 428614
rect 382542 428378 382574 428614
rect 381954 428294 382574 428378
rect 381954 428058 381986 428294
rect 382222 428058 382306 428294
rect 382542 428058 382574 428294
rect 381954 392614 382574 428058
rect 381954 392378 381986 392614
rect 382222 392378 382306 392614
rect 382542 392378 382574 392614
rect 381954 392294 382574 392378
rect 381954 392058 381986 392294
rect 382222 392058 382306 392294
rect 382542 392058 382574 392294
rect 381954 356614 382574 392058
rect 381954 356378 381986 356614
rect 382222 356378 382306 356614
rect 382542 356378 382574 356614
rect 381954 356294 382574 356378
rect 381954 356058 381986 356294
rect 382222 356058 382306 356294
rect 382542 356058 382574 356294
rect 381954 320614 382574 356058
rect 381954 320378 381986 320614
rect 382222 320378 382306 320614
rect 382542 320378 382574 320614
rect 381954 320294 382574 320378
rect 381954 320058 381986 320294
rect 382222 320058 382306 320294
rect 382542 320058 382574 320294
rect 381954 284614 382574 320058
rect 381954 284378 381986 284614
rect 382222 284378 382306 284614
rect 382542 284378 382574 284614
rect 381954 284294 382574 284378
rect 381954 284058 381986 284294
rect 382222 284058 382306 284294
rect 382542 284058 382574 284294
rect 381954 248614 382574 284058
rect 381954 248378 381986 248614
rect 382222 248378 382306 248614
rect 382542 248378 382574 248614
rect 381954 248294 382574 248378
rect 381954 248058 381986 248294
rect 382222 248058 382306 248294
rect 382542 248058 382574 248294
rect 381954 212614 382574 248058
rect 381954 212378 381986 212614
rect 382222 212378 382306 212614
rect 382542 212378 382574 212614
rect 381954 212294 382574 212378
rect 381954 212058 381986 212294
rect 382222 212058 382306 212294
rect 382542 212058 382574 212294
rect 381954 176614 382574 212058
rect 381954 176378 381986 176614
rect 382222 176378 382306 176614
rect 382542 176378 382574 176614
rect 381954 176294 382574 176378
rect 381954 176058 381986 176294
rect 382222 176058 382306 176294
rect 382542 176058 382574 176294
rect 381954 140614 382574 176058
rect 381954 140378 381986 140614
rect 382222 140378 382306 140614
rect 382542 140378 382574 140614
rect 381954 140294 382574 140378
rect 381954 140058 381986 140294
rect 382222 140058 382306 140294
rect 382542 140058 382574 140294
rect 381954 104614 382574 140058
rect 381954 104378 381986 104614
rect 382222 104378 382306 104614
rect 382542 104378 382574 104614
rect 381954 104294 382574 104378
rect 381954 104058 381986 104294
rect 382222 104058 382306 104294
rect 382542 104058 382574 104294
rect 381954 68614 382574 104058
rect 381954 68378 381986 68614
rect 382222 68378 382306 68614
rect 382542 68378 382574 68614
rect 381954 68294 382574 68378
rect 381954 68058 381986 68294
rect 382222 68058 382306 68294
rect 382542 68058 382574 68294
rect 381954 32614 382574 68058
rect 381954 32378 381986 32614
rect 382222 32378 382306 32614
rect 382542 32378 382574 32614
rect 381954 32294 382574 32378
rect 381954 32058 381986 32294
rect 382222 32058 382306 32294
rect 382542 32058 382574 32294
rect 378234 -5382 378266 -5146
rect 378502 -5382 378586 -5146
rect 378822 -5382 378854 -5146
rect 378234 -5466 378854 -5382
rect 378234 -5702 378266 -5466
rect 378502 -5702 378586 -5466
rect 378822 -5702 378854 -5466
rect 378234 -5734 378854 -5702
rect 371954 -6342 371986 -6106
rect 372222 -6342 372306 -6106
rect 372542 -6342 372574 -6106
rect 371954 -6426 372574 -6342
rect 371954 -6662 371986 -6426
rect 372222 -6662 372306 -6426
rect 372542 -6662 372574 -6426
rect 371954 -7654 372574 -6662
rect 381954 -7066 382574 32058
rect 384514 706758 385134 707750
rect 384514 706522 384546 706758
rect 384782 706522 384866 706758
rect 385102 706522 385134 706758
rect 384514 706438 385134 706522
rect 384514 706202 384546 706438
rect 384782 706202 384866 706438
rect 385102 706202 385134 706438
rect 384514 691174 385134 706202
rect 384514 690938 384546 691174
rect 384782 690938 384866 691174
rect 385102 690938 385134 691174
rect 384514 690854 385134 690938
rect 384514 690618 384546 690854
rect 384782 690618 384866 690854
rect 385102 690618 385134 690854
rect 384514 655174 385134 690618
rect 384514 654938 384546 655174
rect 384782 654938 384866 655174
rect 385102 654938 385134 655174
rect 384514 654854 385134 654938
rect 384514 654618 384546 654854
rect 384782 654618 384866 654854
rect 385102 654618 385134 654854
rect 384514 619174 385134 654618
rect 384514 618938 384546 619174
rect 384782 618938 384866 619174
rect 385102 618938 385134 619174
rect 384514 618854 385134 618938
rect 384514 618618 384546 618854
rect 384782 618618 384866 618854
rect 385102 618618 385134 618854
rect 384514 583174 385134 618618
rect 384514 582938 384546 583174
rect 384782 582938 384866 583174
rect 385102 582938 385134 583174
rect 384514 582854 385134 582938
rect 384514 582618 384546 582854
rect 384782 582618 384866 582854
rect 385102 582618 385134 582854
rect 384514 547174 385134 582618
rect 384514 546938 384546 547174
rect 384782 546938 384866 547174
rect 385102 546938 385134 547174
rect 384514 546854 385134 546938
rect 384514 546618 384546 546854
rect 384782 546618 384866 546854
rect 385102 546618 385134 546854
rect 384514 511174 385134 546618
rect 384514 510938 384546 511174
rect 384782 510938 384866 511174
rect 385102 510938 385134 511174
rect 384514 510854 385134 510938
rect 384514 510618 384546 510854
rect 384782 510618 384866 510854
rect 385102 510618 385134 510854
rect 384514 475174 385134 510618
rect 384514 474938 384546 475174
rect 384782 474938 384866 475174
rect 385102 474938 385134 475174
rect 384514 474854 385134 474938
rect 384514 474618 384546 474854
rect 384782 474618 384866 474854
rect 385102 474618 385134 474854
rect 384514 439174 385134 474618
rect 384514 438938 384546 439174
rect 384782 438938 384866 439174
rect 385102 438938 385134 439174
rect 384514 438854 385134 438938
rect 384514 438618 384546 438854
rect 384782 438618 384866 438854
rect 385102 438618 385134 438854
rect 384514 403174 385134 438618
rect 384514 402938 384546 403174
rect 384782 402938 384866 403174
rect 385102 402938 385134 403174
rect 384514 402854 385134 402938
rect 384514 402618 384546 402854
rect 384782 402618 384866 402854
rect 385102 402618 385134 402854
rect 384514 367174 385134 402618
rect 384514 366938 384546 367174
rect 384782 366938 384866 367174
rect 385102 366938 385134 367174
rect 384514 366854 385134 366938
rect 384514 366618 384546 366854
rect 384782 366618 384866 366854
rect 385102 366618 385134 366854
rect 384514 331174 385134 366618
rect 384514 330938 384546 331174
rect 384782 330938 384866 331174
rect 385102 330938 385134 331174
rect 384514 330854 385134 330938
rect 384514 330618 384546 330854
rect 384782 330618 384866 330854
rect 385102 330618 385134 330854
rect 384514 295174 385134 330618
rect 384514 294938 384546 295174
rect 384782 294938 384866 295174
rect 385102 294938 385134 295174
rect 384514 294854 385134 294938
rect 384514 294618 384546 294854
rect 384782 294618 384866 294854
rect 385102 294618 385134 294854
rect 384514 259174 385134 294618
rect 384514 258938 384546 259174
rect 384782 258938 384866 259174
rect 385102 258938 385134 259174
rect 384514 258854 385134 258938
rect 384514 258618 384546 258854
rect 384782 258618 384866 258854
rect 385102 258618 385134 258854
rect 384514 223174 385134 258618
rect 384514 222938 384546 223174
rect 384782 222938 384866 223174
rect 385102 222938 385134 223174
rect 384514 222854 385134 222938
rect 384514 222618 384546 222854
rect 384782 222618 384866 222854
rect 385102 222618 385134 222854
rect 384514 187174 385134 222618
rect 384514 186938 384546 187174
rect 384782 186938 384866 187174
rect 385102 186938 385134 187174
rect 384514 186854 385134 186938
rect 384514 186618 384546 186854
rect 384782 186618 384866 186854
rect 385102 186618 385134 186854
rect 384514 151174 385134 186618
rect 384514 150938 384546 151174
rect 384782 150938 384866 151174
rect 385102 150938 385134 151174
rect 384514 150854 385134 150938
rect 384514 150618 384546 150854
rect 384782 150618 384866 150854
rect 385102 150618 385134 150854
rect 384514 115174 385134 150618
rect 384514 114938 384546 115174
rect 384782 114938 384866 115174
rect 385102 114938 385134 115174
rect 384514 114854 385134 114938
rect 384514 114618 384546 114854
rect 384782 114618 384866 114854
rect 385102 114618 385134 114854
rect 384514 79174 385134 114618
rect 384514 78938 384546 79174
rect 384782 78938 384866 79174
rect 385102 78938 385134 79174
rect 384514 78854 385134 78938
rect 384514 78618 384546 78854
rect 384782 78618 384866 78854
rect 385102 78618 385134 78854
rect 384514 43174 385134 78618
rect 384514 42938 384546 43174
rect 384782 42938 384866 43174
rect 385102 42938 385134 43174
rect 384514 42854 385134 42938
rect 384514 42618 384546 42854
rect 384782 42618 384866 42854
rect 385102 42618 385134 42854
rect 384514 7174 385134 42618
rect 384514 6938 384546 7174
rect 384782 6938 384866 7174
rect 385102 6938 385134 7174
rect 384514 6854 385134 6938
rect 384514 6618 384546 6854
rect 384782 6618 384866 6854
rect 385102 6618 385134 6854
rect 384514 -2266 385134 6618
rect 384514 -2502 384546 -2266
rect 384782 -2502 384866 -2266
rect 385102 -2502 385134 -2266
rect 384514 -2586 385134 -2502
rect 384514 -2822 384546 -2586
rect 384782 -2822 384866 -2586
rect 385102 -2822 385134 -2586
rect 384514 -3814 385134 -2822
rect 388234 694894 388854 708122
rect 388234 694658 388266 694894
rect 388502 694658 388586 694894
rect 388822 694658 388854 694894
rect 388234 694574 388854 694658
rect 388234 694338 388266 694574
rect 388502 694338 388586 694574
rect 388822 694338 388854 694574
rect 388234 658894 388854 694338
rect 388234 658658 388266 658894
rect 388502 658658 388586 658894
rect 388822 658658 388854 658894
rect 388234 658574 388854 658658
rect 388234 658338 388266 658574
rect 388502 658338 388586 658574
rect 388822 658338 388854 658574
rect 388234 622894 388854 658338
rect 388234 622658 388266 622894
rect 388502 622658 388586 622894
rect 388822 622658 388854 622894
rect 388234 622574 388854 622658
rect 388234 622338 388266 622574
rect 388502 622338 388586 622574
rect 388822 622338 388854 622574
rect 388234 586894 388854 622338
rect 388234 586658 388266 586894
rect 388502 586658 388586 586894
rect 388822 586658 388854 586894
rect 388234 586574 388854 586658
rect 388234 586338 388266 586574
rect 388502 586338 388586 586574
rect 388822 586338 388854 586574
rect 388234 550894 388854 586338
rect 388234 550658 388266 550894
rect 388502 550658 388586 550894
rect 388822 550658 388854 550894
rect 388234 550574 388854 550658
rect 388234 550338 388266 550574
rect 388502 550338 388586 550574
rect 388822 550338 388854 550574
rect 388234 514894 388854 550338
rect 388234 514658 388266 514894
rect 388502 514658 388586 514894
rect 388822 514658 388854 514894
rect 388234 514574 388854 514658
rect 388234 514338 388266 514574
rect 388502 514338 388586 514574
rect 388822 514338 388854 514574
rect 388234 478894 388854 514338
rect 388234 478658 388266 478894
rect 388502 478658 388586 478894
rect 388822 478658 388854 478894
rect 388234 478574 388854 478658
rect 388234 478338 388266 478574
rect 388502 478338 388586 478574
rect 388822 478338 388854 478574
rect 388234 442894 388854 478338
rect 388234 442658 388266 442894
rect 388502 442658 388586 442894
rect 388822 442658 388854 442894
rect 388234 442574 388854 442658
rect 388234 442338 388266 442574
rect 388502 442338 388586 442574
rect 388822 442338 388854 442574
rect 388234 406894 388854 442338
rect 388234 406658 388266 406894
rect 388502 406658 388586 406894
rect 388822 406658 388854 406894
rect 388234 406574 388854 406658
rect 388234 406338 388266 406574
rect 388502 406338 388586 406574
rect 388822 406338 388854 406574
rect 388234 370894 388854 406338
rect 388234 370658 388266 370894
rect 388502 370658 388586 370894
rect 388822 370658 388854 370894
rect 388234 370574 388854 370658
rect 388234 370338 388266 370574
rect 388502 370338 388586 370574
rect 388822 370338 388854 370574
rect 388234 334894 388854 370338
rect 388234 334658 388266 334894
rect 388502 334658 388586 334894
rect 388822 334658 388854 334894
rect 388234 334574 388854 334658
rect 388234 334338 388266 334574
rect 388502 334338 388586 334574
rect 388822 334338 388854 334574
rect 388234 298894 388854 334338
rect 388234 298658 388266 298894
rect 388502 298658 388586 298894
rect 388822 298658 388854 298894
rect 388234 298574 388854 298658
rect 388234 298338 388266 298574
rect 388502 298338 388586 298574
rect 388822 298338 388854 298574
rect 388234 262894 388854 298338
rect 388234 262658 388266 262894
rect 388502 262658 388586 262894
rect 388822 262658 388854 262894
rect 388234 262574 388854 262658
rect 388234 262338 388266 262574
rect 388502 262338 388586 262574
rect 388822 262338 388854 262574
rect 388234 226894 388854 262338
rect 388234 226658 388266 226894
rect 388502 226658 388586 226894
rect 388822 226658 388854 226894
rect 388234 226574 388854 226658
rect 388234 226338 388266 226574
rect 388502 226338 388586 226574
rect 388822 226338 388854 226574
rect 388234 190894 388854 226338
rect 388234 190658 388266 190894
rect 388502 190658 388586 190894
rect 388822 190658 388854 190894
rect 388234 190574 388854 190658
rect 388234 190338 388266 190574
rect 388502 190338 388586 190574
rect 388822 190338 388854 190574
rect 388234 154894 388854 190338
rect 388234 154658 388266 154894
rect 388502 154658 388586 154894
rect 388822 154658 388854 154894
rect 388234 154574 388854 154658
rect 388234 154338 388266 154574
rect 388502 154338 388586 154574
rect 388822 154338 388854 154574
rect 388234 118894 388854 154338
rect 388234 118658 388266 118894
rect 388502 118658 388586 118894
rect 388822 118658 388854 118894
rect 388234 118574 388854 118658
rect 388234 118338 388266 118574
rect 388502 118338 388586 118574
rect 388822 118338 388854 118574
rect 388234 82894 388854 118338
rect 388234 82658 388266 82894
rect 388502 82658 388586 82894
rect 388822 82658 388854 82894
rect 388234 82574 388854 82658
rect 388234 82338 388266 82574
rect 388502 82338 388586 82574
rect 388822 82338 388854 82574
rect 388234 46894 388854 82338
rect 388234 46658 388266 46894
rect 388502 46658 388586 46894
rect 388822 46658 388854 46894
rect 388234 46574 388854 46658
rect 388234 46338 388266 46574
rect 388502 46338 388586 46574
rect 388822 46338 388854 46574
rect 388234 10894 388854 46338
rect 388234 10658 388266 10894
rect 388502 10658 388586 10894
rect 388822 10658 388854 10894
rect 388234 10574 388854 10658
rect 388234 10338 388266 10574
rect 388502 10338 388586 10574
rect 388822 10338 388854 10574
rect 388234 -4186 388854 10338
rect 390794 705798 391414 705830
rect 390794 705562 390826 705798
rect 391062 705562 391146 705798
rect 391382 705562 391414 705798
rect 390794 705478 391414 705562
rect 390794 705242 390826 705478
rect 391062 705242 391146 705478
rect 391382 705242 391414 705478
rect 390794 669454 391414 705242
rect 390794 669218 390826 669454
rect 391062 669218 391146 669454
rect 391382 669218 391414 669454
rect 390794 669134 391414 669218
rect 390794 668898 390826 669134
rect 391062 668898 391146 669134
rect 391382 668898 391414 669134
rect 390794 633454 391414 668898
rect 390794 633218 390826 633454
rect 391062 633218 391146 633454
rect 391382 633218 391414 633454
rect 390794 633134 391414 633218
rect 390794 632898 390826 633134
rect 391062 632898 391146 633134
rect 391382 632898 391414 633134
rect 390794 597454 391414 632898
rect 390794 597218 390826 597454
rect 391062 597218 391146 597454
rect 391382 597218 391414 597454
rect 390794 597134 391414 597218
rect 390794 596898 390826 597134
rect 391062 596898 391146 597134
rect 391382 596898 391414 597134
rect 390794 561454 391414 596898
rect 390794 561218 390826 561454
rect 391062 561218 391146 561454
rect 391382 561218 391414 561454
rect 390794 561134 391414 561218
rect 390794 560898 390826 561134
rect 391062 560898 391146 561134
rect 391382 560898 391414 561134
rect 390794 525454 391414 560898
rect 390794 525218 390826 525454
rect 391062 525218 391146 525454
rect 391382 525218 391414 525454
rect 390794 525134 391414 525218
rect 390794 524898 390826 525134
rect 391062 524898 391146 525134
rect 391382 524898 391414 525134
rect 390794 489454 391414 524898
rect 390794 489218 390826 489454
rect 391062 489218 391146 489454
rect 391382 489218 391414 489454
rect 390794 489134 391414 489218
rect 390794 488898 390826 489134
rect 391062 488898 391146 489134
rect 391382 488898 391414 489134
rect 390794 453454 391414 488898
rect 390794 453218 390826 453454
rect 391062 453218 391146 453454
rect 391382 453218 391414 453454
rect 390794 453134 391414 453218
rect 390794 452898 390826 453134
rect 391062 452898 391146 453134
rect 391382 452898 391414 453134
rect 390794 417454 391414 452898
rect 390794 417218 390826 417454
rect 391062 417218 391146 417454
rect 391382 417218 391414 417454
rect 390794 417134 391414 417218
rect 390794 416898 390826 417134
rect 391062 416898 391146 417134
rect 391382 416898 391414 417134
rect 390794 381454 391414 416898
rect 390794 381218 390826 381454
rect 391062 381218 391146 381454
rect 391382 381218 391414 381454
rect 390794 381134 391414 381218
rect 390794 380898 390826 381134
rect 391062 380898 391146 381134
rect 391382 380898 391414 381134
rect 390794 345454 391414 380898
rect 390794 345218 390826 345454
rect 391062 345218 391146 345454
rect 391382 345218 391414 345454
rect 390794 345134 391414 345218
rect 390794 344898 390826 345134
rect 391062 344898 391146 345134
rect 391382 344898 391414 345134
rect 390794 309454 391414 344898
rect 390794 309218 390826 309454
rect 391062 309218 391146 309454
rect 391382 309218 391414 309454
rect 390794 309134 391414 309218
rect 390794 308898 390826 309134
rect 391062 308898 391146 309134
rect 391382 308898 391414 309134
rect 390794 273454 391414 308898
rect 390794 273218 390826 273454
rect 391062 273218 391146 273454
rect 391382 273218 391414 273454
rect 390794 273134 391414 273218
rect 390794 272898 390826 273134
rect 391062 272898 391146 273134
rect 391382 272898 391414 273134
rect 390794 237454 391414 272898
rect 390794 237218 390826 237454
rect 391062 237218 391146 237454
rect 391382 237218 391414 237454
rect 390794 237134 391414 237218
rect 390794 236898 390826 237134
rect 391062 236898 391146 237134
rect 391382 236898 391414 237134
rect 390794 201454 391414 236898
rect 390794 201218 390826 201454
rect 391062 201218 391146 201454
rect 391382 201218 391414 201454
rect 390794 201134 391414 201218
rect 390794 200898 390826 201134
rect 391062 200898 391146 201134
rect 391382 200898 391414 201134
rect 390794 165454 391414 200898
rect 390794 165218 390826 165454
rect 391062 165218 391146 165454
rect 391382 165218 391414 165454
rect 390794 165134 391414 165218
rect 390794 164898 390826 165134
rect 391062 164898 391146 165134
rect 391382 164898 391414 165134
rect 390794 129454 391414 164898
rect 390794 129218 390826 129454
rect 391062 129218 391146 129454
rect 391382 129218 391414 129454
rect 390794 129134 391414 129218
rect 390794 128898 390826 129134
rect 391062 128898 391146 129134
rect 391382 128898 391414 129134
rect 390794 93454 391414 128898
rect 390794 93218 390826 93454
rect 391062 93218 391146 93454
rect 391382 93218 391414 93454
rect 390794 93134 391414 93218
rect 390794 92898 390826 93134
rect 391062 92898 391146 93134
rect 391382 92898 391414 93134
rect 390794 57454 391414 92898
rect 390794 57218 390826 57454
rect 391062 57218 391146 57454
rect 391382 57218 391414 57454
rect 390794 57134 391414 57218
rect 390794 56898 390826 57134
rect 391062 56898 391146 57134
rect 391382 56898 391414 57134
rect 390794 21454 391414 56898
rect 390794 21218 390826 21454
rect 391062 21218 391146 21454
rect 391382 21218 391414 21454
rect 390794 21134 391414 21218
rect 390794 20898 390826 21134
rect 391062 20898 391146 21134
rect 391382 20898 391414 21134
rect 390794 -1306 391414 20898
rect 390794 -1542 390826 -1306
rect 391062 -1542 391146 -1306
rect 391382 -1542 391414 -1306
rect 390794 -1626 391414 -1542
rect 390794 -1862 390826 -1626
rect 391062 -1862 391146 -1626
rect 391382 -1862 391414 -1626
rect 390794 -1894 391414 -1862
rect 391954 698614 392574 710042
rect 401954 711558 402574 711590
rect 401954 711322 401986 711558
rect 402222 711322 402306 711558
rect 402542 711322 402574 711558
rect 401954 711238 402574 711322
rect 401954 711002 401986 711238
rect 402222 711002 402306 711238
rect 402542 711002 402574 711238
rect 398234 709638 398854 709670
rect 398234 709402 398266 709638
rect 398502 709402 398586 709638
rect 398822 709402 398854 709638
rect 398234 709318 398854 709402
rect 398234 709082 398266 709318
rect 398502 709082 398586 709318
rect 398822 709082 398854 709318
rect 391954 698378 391986 698614
rect 392222 698378 392306 698614
rect 392542 698378 392574 698614
rect 391954 698294 392574 698378
rect 391954 698058 391986 698294
rect 392222 698058 392306 698294
rect 392542 698058 392574 698294
rect 391954 662614 392574 698058
rect 391954 662378 391986 662614
rect 392222 662378 392306 662614
rect 392542 662378 392574 662614
rect 391954 662294 392574 662378
rect 391954 662058 391986 662294
rect 392222 662058 392306 662294
rect 392542 662058 392574 662294
rect 391954 626614 392574 662058
rect 391954 626378 391986 626614
rect 392222 626378 392306 626614
rect 392542 626378 392574 626614
rect 391954 626294 392574 626378
rect 391954 626058 391986 626294
rect 392222 626058 392306 626294
rect 392542 626058 392574 626294
rect 391954 590614 392574 626058
rect 391954 590378 391986 590614
rect 392222 590378 392306 590614
rect 392542 590378 392574 590614
rect 391954 590294 392574 590378
rect 391954 590058 391986 590294
rect 392222 590058 392306 590294
rect 392542 590058 392574 590294
rect 391954 554614 392574 590058
rect 391954 554378 391986 554614
rect 392222 554378 392306 554614
rect 392542 554378 392574 554614
rect 391954 554294 392574 554378
rect 391954 554058 391986 554294
rect 392222 554058 392306 554294
rect 392542 554058 392574 554294
rect 391954 518614 392574 554058
rect 391954 518378 391986 518614
rect 392222 518378 392306 518614
rect 392542 518378 392574 518614
rect 391954 518294 392574 518378
rect 391954 518058 391986 518294
rect 392222 518058 392306 518294
rect 392542 518058 392574 518294
rect 391954 482614 392574 518058
rect 391954 482378 391986 482614
rect 392222 482378 392306 482614
rect 392542 482378 392574 482614
rect 391954 482294 392574 482378
rect 391954 482058 391986 482294
rect 392222 482058 392306 482294
rect 392542 482058 392574 482294
rect 391954 446614 392574 482058
rect 391954 446378 391986 446614
rect 392222 446378 392306 446614
rect 392542 446378 392574 446614
rect 391954 446294 392574 446378
rect 391954 446058 391986 446294
rect 392222 446058 392306 446294
rect 392542 446058 392574 446294
rect 391954 410614 392574 446058
rect 391954 410378 391986 410614
rect 392222 410378 392306 410614
rect 392542 410378 392574 410614
rect 391954 410294 392574 410378
rect 391954 410058 391986 410294
rect 392222 410058 392306 410294
rect 392542 410058 392574 410294
rect 391954 374614 392574 410058
rect 391954 374378 391986 374614
rect 392222 374378 392306 374614
rect 392542 374378 392574 374614
rect 391954 374294 392574 374378
rect 391954 374058 391986 374294
rect 392222 374058 392306 374294
rect 392542 374058 392574 374294
rect 391954 338614 392574 374058
rect 391954 338378 391986 338614
rect 392222 338378 392306 338614
rect 392542 338378 392574 338614
rect 391954 338294 392574 338378
rect 391954 338058 391986 338294
rect 392222 338058 392306 338294
rect 392542 338058 392574 338294
rect 391954 302614 392574 338058
rect 391954 302378 391986 302614
rect 392222 302378 392306 302614
rect 392542 302378 392574 302614
rect 391954 302294 392574 302378
rect 391954 302058 391986 302294
rect 392222 302058 392306 302294
rect 392542 302058 392574 302294
rect 391954 266614 392574 302058
rect 391954 266378 391986 266614
rect 392222 266378 392306 266614
rect 392542 266378 392574 266614
rect 391954 266294 392574 266378
rect 391954 266058 391986 266294
rect 392222 266058 392306 266294
rect 392542 266058 392574 266294
rect 391954 230614 392574 266058
rect 391954 230378 391986 230614
rect 392222 230378 392306 230614
rect 392542 230378 392574 230614
rect 391954 230294 392574 230378
rect 391954 230058 391986 230294
rect 392222 230058 392306 230294
rect 392542 230058 392574 230294
rect 391954 194614 392574 230058
rect 391954 194378 391986 194614
rect 392222 194378 392306 194614
rect 392542 194378 392574 194614
rect 391954 194294 392574 194378
rect 391954 194058 391986 194294
rect 392222 194058 392306 194294
rect 392542 194058 392574 194294
rect 391954 158614 392574 194058
rect 391954 158378 391986 158614
rect 392222 158378 392306 158614
rect 392542 158378 392574 158614
rect 391954 158294 392574 158378
rect 391954 158058 391986 158294
rect 392222 158058 392306 158294
rect 392542 158058 392574 158294
rect 391954 122614 392574 158058
rect 391954 122378 391986 122614
rect 392222 122378 392306 122614
rect 392542 122378 392574 122614
rect 391954 122294 392574 122378
rect 391954 122058 391986 122294
rect 392222 122058 392306 122294
rect 392542 122058 392574 122294
rect 391954 86614 392574 122058
rect 391954 86378 391986 86614
rect 392222 86378 392306 86614
rect 392542 86378 392574 86614
rect 391954 86294 392574 86378
rect 391954 86058 391986 86294
rect 392222 86058 392306 86294
rect 392542 86058 392574 86294
rect 391954 50614 392574 86058
rect 391954 50378 391986 50614
rect 392222 50378 392306 50614
rect 392542 50378 392574 50614
rect 391954 50294 392574 50378
rect 391954 50058 391986 50294
rect 392222 50058 392306 50294
rect 392542 50058 392574 50294
rect 391954 14614 392574 50058
rect 391954 14378 391986 14614
rect 392222 14378 392306 14614
rect 392542 14378 392574 14614
rect 391954 14294 392574 14378
rect 391954 14058 391986 14294
rect 392222 14058 392306 14294
rect 392542 14058 392574 14294
rect 388234 -4422 388266 -4186
rect 388502 -4422 388586 -4186
rect 388822 -4422 388854 -4186
rect 388234 -4506 388854 -4422
rect 388234 -4742 388266 -4506
rect 388502 -4742 388586 -4506
rect 388822 -4742 388854 -4506
rect 388234 -5734 388854 -4742
rect 381954 -7302 381986 -7066
rect 382222 -7302 382306 -7066
rect 382542 -7302 382574 -7066
rect 381954 -7386 382574 -7302
rect 381954 -7622 381986 -7386
rect 382222 -7622 382306 -7386
rect 382542 -7622 382574 -7386
rect 381954 -7654 382574 -7622
rect 391954 -6106 392574 14058
rect 394514 707718 395134 707750
rect 394514 707482 394546 707718
rect 394782 707482 394866 707718
rect 395102 707482 395134 707718
rect 394514 707398 395134 707482
rect 394514 707162 394546 707398
rect 394782 707162 394866 707398
rect 395102 707162 395134 707398
rect 394514 673174 395134 707162
rect 394514 672938 394546 673174
rect 394782 672938 394866 673174
rect 395102 672938 395134 673174
rect 394514 672854 395134 672938
rect 394514 672618 394546 672854
rect 394782 672618 394866 672854
rect 395102 672618 395134 672854
rect 394514 637174 395134 672618
rect 394514 636938 394546 637174
rect 394782 636938 394866 637174
rect 395102 636938 395134 637174
rect 394514 636854 395134 636938
rect 394514 636618 394546 636854
rect 394782 636618 394866 636854
rect 395102 636618 395134 636854
rect 394514 601174 395134 636618
rect 394514 600938 394546 601174
rect 394782 600938 394866 601174
rect 395102 600938 395134 601174
rect 394514 600854 395134 600938
rect 394514 600618 394546 600854
rect 394782 600618 394866 600854
rect 395102 600618 395134 600854
rect 394514 565174 395134 600618
rect 394514 564938 394546 565174
rect 394782 564938 394866 565174
rect 395102 564938 395134 565174
rect 394514 564854 395134 564938
rect 394514 564618 394546 564854
rect 394782 564618 394866 564854
rect 395102 564618 395134 564854
rect 394514 529174 395134 564618
rect 394514 528938 394546 529174
rect 394782 528938 394866 529174
rect 395102 528938 395134 529174
rect 394514 528854 395134 528938
rect 394514 528618 394546 528854
rect 394782 528618 394866 528854
rect 395102 528618 395134 528854
rect 394514 493174 395134 528618
rect 394514 492938 394546 493174
rect 394782 492938 394866 493174
rect 395102 492938 395134 493174
rect 394514 492854 395134 492938
rect 394514 492618 394546 492854
rect 394782 492618 394866 492854
rect 395102 492618 395134 492854
rect 394514 457174 395134 492618
rect 394514 456938 394546 457174
rect 394782 456938 394866 457174
rect 395102 456938 395134 457174
rect 394514 456854 395134 456938
rect 394514 456618 394546 456854
rect 394782 456618 394866 456854
rect 395102 456618 395134 456854
rect 394514 421174 395134 456618
rect 394514 420938 394546 421174
rect 394782 420938 394866 421174
rect 395102 420938 395134 421174
rect 394514 420854 395134 420938
rect 394514 420618 394546 420854
rect 394782 420618 394866 420854
rect 395102 420618 395134 420854
rect 394514 385174 395134 420618
rect 394514 384938 394546 385174
rect 394782 384938 394866 385174
rect 395102 384938 395134 385174
rect 394514 384854 395134 384938
rect 394514 384618 394546 384854
rect 394782 384618 394866 384854
rect 395102 384618 395134 384854
rect 394514 349174 395134 384618
rect 394514 348938 394546 349174
rect 394782 348938 394866 349174
rect 395102 348938 395134 349174
rect 394514 348854 395134 348938
rect 394514 348618 394546 348854
rect 394782 348618 394866 348854
rect 395102 348618 395134 348854
rect 394514 313174 395134 348618
rect 394514 312938 394546 313174
rect 394782 312938 394866 313174
rect 395102 312938 395134 313174
rect 394514 312854 395134 312938
rect 394514 312618 394546 312854
rect 394782 312618 394866 312854
rect 395102 312618 395134 312854
rect 394514 277174 395134 312618
rect 394514 276938 394546 277174
rect 394782 276938 394866 277174
rect 395102 276938 395134 277174
rect 394514 276854 395134 276938
rect 394514 276618 394546 276854
rect 394782 276618 394866 276854
rect 395102 276618 395134 276854
rect 394514 241174 395134 276618
rect 394514 240938 394546 241174
rect 394782 240938 394866 241174
rect 395102 240938 395134 241174
rect 394514 240854 395134 240938
rect 394514 240618 394546 240854
rect 394782 240618 394866 240854
rect 395102 240618 395134 240854
rect 394514 205174 395134 240618
rect 394514 204938 394546 205174
rect 394782 204938 394866 205174
rect 395102 204938 395134 205174
rect 394514 204854 395134 204938
rect 394514 204618 394546 204854
rect 394782 204618 394866 204854
rect 395102 204618 395134 204854
rect 394514 169174 395134 204618
rect 394514 168938 394546 169174
rect 394782 168938 394866 169174
rect 395102 168938 395134 169174
rect 394514 168854 395134 168938
rect 394514 168618 394546 168854
rect 394782 168618 394866 168854
rect 395102 168618 395134 168854
rect 394514 133174 395134 168618
rect 394514 132938 394546 133174
rect 394782 132938 394866 133174
rect 395102 132938 395134 133174
rect 394514 132854 395134 132938
rect 394514 132618 394546 132854
rect 394782 132618 394866 132854
rect 395102 132618 395134 132854
rect 394514 97174 395134 132618
rect 394514 96938 394546 97174
rect 394782 96938 394866 97174
rect 395102 96938 395134 97174
rect 394514 96854 395134 96938
rect 394514 96618 394546 96854
rect 394782 96618 394866 96854
rect 395102 96618 395134 96854
rect 394514 61174 395134 96618
rect 394514 60938 394546 61174
rect 394782 60938 394866 61174
rect 395102 60938 395134 61174
rect 394514 60854 395134 60938
rect 394514 60618 394546 60854
rect 394782 60618 394866 60854
rect 395102 60618 395134 60854
rect 394514 25174 395134 60618
rect 394514 24938 394546 25174
rect 394782 24938 394866 25174
rect 395102 24938 395134 25174
rect 394514 24854 395134 24938
rect 394514 24618 394546 24854
rect 394782 24618 394866 24854
rect 395102 24618 395134 24854
rect 394514 -3226 395134 24618
rect 394514 -3462 394546 -3226
rect 394782 -3462 394866 -3226
rect 395102 -3462 395134 -3226
rect 394514 -3546 395134 -3462
rect 394514 -3782 394546 -3546
rect 394782 -3782 394866 -3546
rect 395102 -3782 395134 -3546
rect 394514 -3814 395134 -3782
rect 398234 676894 398854 709082
rect 398234 676658 398266 676894
rect 398502 676658 398586 676894
rect 398822 676658 398854 676894
rect 398234 676574 398854 676658
rect 398234 676338 398266 676574
rect 398502 676338 398586 676574
rect 398822 676338 398854 676574
rect 398234 640894 398854 676338
rect 398234 640658 398266 640894
rect 398502 640658 398586 640894
rect 398822 640658 398854 640894
rect 398234 640574 398854 640658
rect 398234 640338 398266 640574
rect 398502 640338 398586 640574
rect 398822 640338 398854 640574
rect 398234 604894 398854 640338
rect 398234 604658 398266 604894
rect 398502 604658 398586 604894
rect 398822 604658 398854 604894
rect 398234 604574 398854 604658
rect 398234 604338 398266 604574
rect 398502 604338 398586 604574
rect 398822 604338 398854 604574
rect 398234 568894 398854 604338
rect 398234 568658 398266 568894
rect 398502 568658 398586 568894
rect 398822 568658 398854 568894
rect 398234 568574 398854 568658
rect 398234 568338 398266 568574
rect 398502 568338 398586 568574
rect 398822 568338 398854 568574
rect 398234 532894 398854 568338
rect 398234 532658 398266 532894
rect 398502 532658 398586 532894
rect 398822 532658 398854 532894
rect 398234 532574 398854 532658
rect 398234 532338 398266 532574
rect 398502 532338 398586 532574
rect 398822 532338 398854 532574
rect 398234 496894 398854 532338
rect 398234 496658 398266 496894
rect 398502 496658 398586 496894
rect 398822 496658 398854 496894
rect 398234 496574 398854 496658
rect 398234 496338 398266 496574
rect 398502 496338 398586 496574
rect 398822 496338 398854 496574
rect 398234 460894 398854 496338
rect 398234 460658 398266 460894
rect 398502 460658 398586 460894
rect 398822 460658 398854 460894
rect 398234 460574 398854 460658
rect 398234 460338 398266 460574
rect 398502 460338 398586 460574
rect 398822 460338 398854 460574
rect 398234 424894 398854 460338
rect 398234 424658 398266 424894
rect 398502 424658 398586 424894
rect 398822 424658 398854 424894
rect 398234 424574 398854 424658
rect 398234 424338 398266 424574
rect 398502 424338 398586 424574
rect 398822 424338 398854 424574
rect 398234 388894 398854 424338
rect 398234 388658 398266 388894
rect 398502 388658 398586 388894
rect 398822 388658 398854 388894
rect 398234 388574 398854 388658
rect 398234 388338 398266 388574
rect 398502 388338 398586 388574
rect 398822 388338 398854 388574
rect 398234 352894 398854 388338
rect 398234 352658 398266 352894
rect 398502 352658 398586 352894
rect 398822 352658 398854 352894
rect 398234 352574 398854 352658
rect 398234 352338 398266 352574
rect 398502 352338 398586 352574
rect 398822 352338 398854 352574
rect 398234 316894 398854 352338
rect 398234 316658 398266 316894
rect 398502 316658 398586 316894
rect 398822 316658 398854 316894
rect 398234 316574 398854 316658
rect 398234 316338 398266 316574
rect 398502 316338 398586 316574
rect 398822 316338 398854 316574
rect 398234 280894 398854 316338
rect 398234 280658 398266 280894
rect 398502 280658 398586 280894
rect 398822 280658 398854 280894
rect 398234 280574 398854 280658
rect 398234 280338 398266 280574
rect 398502 280338 398586 280574
rect 398822 280338 398854 280574
rect 398234 244894 398854 280338
rect 398234 244658 398266 244894
rect 398502 244658 398586 244894
rect 398822 244658 398854 244894
rect 398234 244574 398854 244658
rect 398234 244338 398266 244574
rect 398502 244338 398586 244574
rect 398822 244338 398854 244574
rect 398234 208894 398854 244338
rect 398234 208658 398266 208894
rect 398502 208658 398586 208894
rect 398822 208658 398854 208894
rect 398234 208574 398854 208658
rect 398234 208338 398266 208574
rect 398502 208338 398586 208574
rect 398822 208338 398854 208574
rect 398234 172894 398854 208338
rect 398234 172658 398266 172894
rect 398502 172658 398586 172894
rect 398822 172658 398854 172894
rect 398234 172574 398854 172658
rect 398234 172338 398266 172574
rect 398502 172338 398586 172574
rect 398822 172338 398854 172574
rect 398234 136894 398854 172338
rect 398234 136658 398266 136894
rect 398502 136658 398586 136894
rect 398822 136658 398854 136894
rect 398234 136574 398854 136658
rect 398234 136338 398266 136574
rect 398502 136338 398586 136574
rect 398822 136338 398854 136574
rect 398234 100894 398854 136338
rect 398234 100658 398266 100894
rect 398502 100658 398586 100894
rect 398822 100658 398854 100894
rect 398234 100574 398854 100658
rect 398234 100338 398266 100574
rect 398502 100338 398586 100574
rect 398822 100338 398854 100574
rect 398234 64894 398854 100338
rect 398234 64658 398266 64894
rect 398502 64658 398586 64894
rect 398822 64658 398854 64894
rect 398234 64574 398854 64658
rect 398234 64338 398266 64574
rect 398502 64338 398586 64574
rect 398822 64338 398854 64574
rect 398234 28894 398854 64338
rect 398234 28658 398266 28894
rect 398502 28658 398586 28894
rect 398822 28658 398854 28894
rect 398234 28574 398854 28658
rect 398234 28338 398266 28574
rect 398502 28338 398586 28574
rect 398822 28338 398854 28574
rect 398234 -5146 398854 28338
rect 400794 704838 401414 705830
rect 400794 704602 400826 704838
rect 401062 704602 401146 704838
rect 401382 704602 401414 704838
rect 400794 704518 401414 704602
rect 400794 704282 400826 704518
rect 401062 704282 401146 704518
rect 401382 704282 401414 704518
rect 400794 687454 401414 704282
rect 400794 687218 400826 687454
rect 401062 687218 401146 687454
rect 401382 687218 401414 687454
rect 400794 687134 401414 687218
rect 400794 686898 400826 687134
rect 401062 686898 401146 687134
rect 401382 686898 401414 687134
rect 400794 651454 401414 686898
rect 400794 651218 400826 651454
rect 401062 651218 401146 651454
rect 401382 651218 401414 651454
rect 400794 651134 401414 651218
rect 400794 650898 400826 651134
rect 401062 650898 401146 651134
rect 401382 650898 401414 651134
rect 400794 615454 401414 650898
rect 400794 615218 400826 615454
rect 401062 615218 401146 615454
rect 401382 615218 401414 615454
rect 400794 615134 401414 615218
rect 400794 614898 400826 615134
rect 401062 614898 401146 615134
rect 401382 614898 401414 615134
rect 400794 579454 401414 614898
rect 400794 579218 400826 579454
rect 401062 579218 401146 579454
rect 401382 579218 401414 579454
rect 400794 579134 401414 579218
rect 400794 578898 400826 579134
rect 401062 578898 401146 579134
rect 401382 578898 401414 579134
rect 400794 543454 401414 578898
rect 400794 543218 400826 543454
rect 401062 543218 401146 543454
rect 401382 543218 401414 543454
rect 400794 543134 401414 543218
rect 400794 542898 400826 543134
rect 401062 542898 401146 543134
rect 401382 542898 401414 543134
rect 400794 507454 401414 542898
rect 400794 507218 400826 507454
rect 401062 507218 401146 507454
rect 401382 507218 401414 507454
rect 400794 507134 401414 507218
rect 400794 506898 400826 507134
rect 401062 506898 401146 507134
rect 401382 506898 401414 507134
rect 400794 471454 401414 506898
rect 400794 471218 400826 471454
rect 401062 471218 401146 471454
rect 401382 471218 401414 471454
rect 400794 471134 401414 471218
rect 400794 470898 400826 471134
rect 401062 470898 401146 471134
rect 401382 470898 401414 471134
rect 400794 435454 401414 470898
rect 400794 435218 400826 435454
rect 401062 435218 401146 435454
rect 401382 435218 401414 435454
rect 400794 435134 401414 435218
rect 400794 434898 400826 435134
rect 401062 434898 401146 435134
rect 401382 434898 401414 435134
rect 400794 399454 401414 434898
rect 400794 399218 400826 399454
rect 401062 399218 401146 399454
rect 401382 399218 401414 399454
rect 400794 399134 401414 399218
rect 400794 398898 400826 399134
rect 401062 398898 401146 399134
rect 401382 398898 401414 399134
rect 400794 363454 401414 398898
rect 400794 363218 400826 363454
rect 401062 363218 401146 363454
rect 401382 363218 401414 363454
rect 400794 363134 401414 363218
rect 400794 362898 400826 363134
rect 401062 362898 401146 363134
rect 401382 362898 401414 363134
rect 400794 327454 401414 362898
rect 400794 327218 400826 327454
rect 401062 327218 401146 327454
rect 401382 327218 401414 327454
rect 400794 327134 401414 327218
rect 400794 326898 400826 327134
rect 401062 326898 401146 327134
rect 401382 326898 401414 327134
rect 400794 291454 401414 326898
rect 400794 291218 400826 291454
rect 401062 291218 401146 291454
rect 401382 291218 401414 291454
rect 400794 291134 401414 291218
rect 400794 290898 400826 291134
rect 401062 290898 401146 291134
rect 401382 290898 401414 291134
rect 400794 255454 401414 290898
rect 400794 255218 400826 255454
rect 401062 255218 401146 255454
rect 401382 255218 401414 255454
rect 400794 255134 401414 255218
rect 400794 254898 400826 255134
rect 401062 254898 401146 255134
rect 401382 254898 401414 255134
rect 400794 219454 401414 254898
rect 400794 219218 400826 219454
rect 401062 219218 401146 219454
rect 401382 219218 401414 219454
rect 400794 219134 401414 219218
rect 400794 218898 400826 219134
rect 401062 218898 401146 219134
rect 401382 218898 401414 219134
rect 400794 183454 401414 218898
rect 400794 183218 400826 183454
rect 401062 183218 401146 183454
rect 401382 183218 401414 183454
rect 400794 183134 401414 183218
rect 400794 182898 400826 183134
rect 401062 182898 401146 183134
rect 401382 182898 401414 183134
rect 400794 147454 401414 182898
rect 400794 147218 400826 147454
rect 401062 147218 401146 147454
rect 401382 147218 401414 147454
rect 400794 147134 401414 147218
rect 400794 146898 400826 147134
rect 401062 146898 401146 147134
rect 401382 146898 401414 147134
rect 400794 111454 401414 146898
rect 400794 111218 400826 111454
rect 401062 111218 401146 111454
rect 401382 111218 401414 111454
rect 400794 111134 401414 111218
rect 400794 110898 400826 111134
rect 401062 110898 401146 111134
rect 401382 110898 401414 111134
rect 400794 75454 401414 110898
rect 400794 75218 400826 75454
rect 401062 75218 401146 75454
rect 401382 75218 401414 75454
rect 400794 75134 401414 75218
rect 400794 74898 400826 75134
rect 401062 74898 401146 75134
rect 401382 74898 401414 75134
rect 400794 39454 401414 74898
rect 400794 39218 400826 39454
rect 401062 39218 401146 39454
rect 401382 39218 401414 39454
rect 400794 39134 401414 39218
rect 400794 38898 400826 39134
rect 401062 38898 401146 39134
rect 401382 38898 401414 39134
rect 400794 3454 401414 38898
rect 400794 3218 400826 3454
rect 401062 3218 401146 3454
rect 401382 3218 401414 3454
rect 400794 3134 401414 3218
rect 400794 2898 400826 3134
rect 401062 2898 401146 3134
rect 401382 2898 401414 3134
rect 400794 -346 401414 2898
rect 400794 -582 400826 -346
rect 401062 -582 401146 -346
rect 401382 -582 401414 -346
rect 400794 -666 401414 -582
rect 400794 -902 400826 -666
rect 401062 -902 401146 -666
rect 401382 -902 401414 -666
rect 400794 -1894 401414 -902
rect 401954 680614 402574 711002
rect 411954 710598 412574 711590
rect 411954 710362 411986 710598
rect 412222 710362 412306 710598
rect 412542 710362 412574 710598
rect 411954 710278 412574 710362
rect 411954 710042 411986 710278
rect 412222 710042 412306 710278
rect 412542 710042 412574 710278
rect 408234 708678 408854 709670
rect 408234 708442 408266 708678
rect 408502 708442 408586 708678
rect 408822 708442 408854 708678
rect 408234 708358 408854 708442
rect 408234 708122 408266 708358
rect 408502 708122 408586 708358
rect 408822 708122 408854 708358
rect 401954 680378 401986 680614
rect 402222 680378 402306 680614
rect 402542 680378 402574 680614
rect 401954 680294 402574 680378
rect 401954 680058 401986 680294
rect 402222 680058 402306 680294
rect 402542 680058 402574 680294
rect 401954 644614 402574 680058
rect 401954 644378 401986 644614
rect 402222 644378 402306 644614
rect 402542 644378 402574 644614
rect 401954 644294 402574 644378
rect 401954 644058 401986 644294
rect 402222 644058 402306 644294
rect 402542 644058 402574 644294
rect 401954 608614 402574 644058
rect 401954 608378 401986 608614
rect 402222 608378 402306 608614
rect 402542 608378 402574 608614
rect 401954 608294 402574 608378
rect 401954 608058 401986 608294
rect 402222 608058 402306 608294
rect 402542 608058 402574 608294
rect 401954 572614 402574 608058
rect 401954 572378 401986 572614
rect 402222 572378 402306 572614
rect 402542 572378 402574 572614
rect 401954 572294 402574 572378
rect 401954 572058 401986 572294
rect 402222 572058 402306 572294
rect 402542 572058 402574 572294
rect 401954 536614 402574 572058
rect 401954 536378 401986 536614
rect 402222 536378 402306 536614
rect 402542 536378 402574 536614
rect 401954 536294 402574 536378
rect 401954 536058 401986 536294
rect 402222 536058 402306 536294
rect 402542 536058 402574 536294
rect 401954 500614 402574 536058
rect 401954 500378 401986 500614
rect 402222 500378 402306 500614
rect 402542 500378 402574 500614
rect 401954 500294 402574 500378
rect 401954 500058 401986 500294
rect 402222 500058 402306 500294
rect 402542 500058 402574 500294
rect 401954 464614 402574 500058
rect 401954 464378 401986 464614
rect 402222 464378 402306 464614
rect 402542 464378 402574 464614
rect 401954 464294 402574 464378
rect 401954 464058 401986 464294
rect 402222 464058 402306 464294
rect 402542 464058 402574 464294
rect 401954 428614 402574 464058
rect 401954 428378 401986 428614
rect 402222 428378 402306 428614
rect 402542 428378 402574 428614
rect 401954 428294 402574 428378
rect 401954 428058 401986 428294
rect 402222 428058 402306 428294
rect 402542 428058 402574 428294
rect 401954 392614 402574 428058
rect 401954 392378 401986 392614
rect 402222 392378 402306 392614
rect 402542 392378 402574 392614
rect 401954 392294 402574 392378
rect 401954 392058 401986 392294
rect 402222 392058 402306 392294
rect 402542 392058 402574 392294
rect 401954 356614 402574 392058
rect 401954 356378 401986 356614
rect 402222 356378 402306 356614
rect 402542 356378 402574 356614
rect 401954 356294 402574 356378
rect 401954 356058 401986 356294
rect 402222 356058 402306 356294
rect 402542 356058 402574 356294
rect 401954 320614 402574 356058
rect 401954 320378 401986 320614
rect 402222 320378 402306 320614
rect 402542 320378 402574 320614
rect 401954 320294 402574 320378
rect 401954 320058 401986 320294
rect 402222 320058 402306 320294
rect 402542 320058 402574 320294
rect 401954 284614 402574 320058
rect 401954 284378 401986 284614
rect 402222 284378 402306 284614
rect 402542 284378 402574 284614
rect 401954 284294 402574 284378
rect 401954 284058 401986 284294
rect 402222 284058 402306 284294
rect 402542 284058 402574 284294
rect 401954 248614 402574 284058
rect 401954 248378 401986 248614
rect 402222 248378 402306 248614
rect 402542 248378 402574 248614
rect 401954 248294 402574 248378
rect 401954 248058 401986 248294
rect 402222 248058 402306 248294
rect 402542 248058 402574 248294
rect 401954 212614 402574 248058
rect 401954 212378 401986 212614
rect 402222 212378 402306 212614
rect 402542 212378 402574 212614
rect 401954 212294 402574 212378
rect 401954 212058 401986 212294
rect 402222 212058 402306 212294
rect 402542 212058 402574 212294
rect 401954 176614 402574 212058
rect 401954 176378 401986 176614
rect 402222 176378 402306 176614
rect 402542 176378 402574 176614
rect 401954 176294 402574 176378
rect 401954 176058 401986 176294
rect 402222 176058 402306 176294
rect 402542 176058 402574 176294
rect 401954 140614 402574 176058
rect 401954 140378 401986 140614
rect 402222 140378 402306 140614
rect 402542 140378 402574 140614
rect 401954 140294 402574 140378
rect 401954 140058 401986 140294
rect 402222 140058 402306 140294
rect 402542 140058 402574 140294
rect 401954 104614 402574 140058
rect 401954 104378 401986 104614
rect 402222 104378 402306 104614
rect 402542 104378 402574 104614
rect 401954 104294 402574 104378
rect 401954 104058 401986 104294
rect 402222 104058 402306 104294
rect 402542 104058 402574 104294
rect 401954 68614 402574 104058
rect 401954 68378 401986 68614
rect 402222 68378 402306 68614
rect 402542 68378 402574 68614
rect 401954 68294 402574 68378
rect 401954 68058 401986 68294
rect 402222 68058 402306 68294
rect 402542 68058 402574 68294
rect 401954 32614 402574 68058
rect 401954 32378 401986 32614
rect 402222 32378 402306 32614
rect 402542 32378 402574 32614
rect 401954 32294 402574 32378
rect 401954 32058 401986 32294
rect 402222 32058 402306 32294
rect 402542 32058 402574 32294
rect 398234 -5382 398266 -5146
rect 398502 -5382 398586 -5146
rect 398822 -5382 398854 -5146
rect 398234 -5466 398854 -5382
rect 398234 -5702 398266 -5466
rect 398502 -5702 398586 -5466
rect 398822 -5702 398854 -5466
rect 398234 -5734 398854 -5702
rect 391954 -6342 391986 -6106
rect 392222 -6342 392306 -6106
rect 392542 -6342 392574 -6106
rect 391954 -6426 392574 -6342
rect 391954 -6662 391986 -6426
rect 392222 -6662 392306 -6426
rect 392542 -6662 392574 -6426
rect 391954 -7654 392574 -6662
rect 401954 -7066 402574 32058
rect 404514 706758 405134 707750
rect 404514 706522 404546 706758
rect 404782 706522 404866 706758
rect 405102 706522 405134 706758
rect 404514 706438 405134 706522
rect 404514 706202 404546 706438
rect 404782 706202 404866 706438
rect 405102 706202 405134 706438
rect 404514 691174 405134 706202
rect 404514 690938 404546 691174
rect 404782 690938 404866 691174
rect 405102 690938 405134 691174
rect 404514 690854 405134 690938
rect 404514 690618 404546 690854
rect 404782 690618 404866 690854
rect 405102 690618 405134 690854
rect 404514 655174 405134 690618
rect 404514 654938 404546 655174
rect 404782 654938 404866 655174
rect 405102 654938 405134 655174
rect 404514 654854 405134 654938
rect 404514 654618 404546 654854
rect 404782 654618 404866 654854
rect 405102 654618 405134 654854
rect 404514 619174 405134 654618
rect 404514 618938 404546 619174
rect 404782 618938 404866 619174
rect 405102 618938 405134 619174
rect 404514 618854 405134 618938
rect 404514 618618 404546 618854
rect 404782 618618 404866 618854
rect 405102 618618 405134 618854
rect 404514 583174 405134 618618
rect 404514 582938 404546 583174
rect 404782 582938 404866 583174
rect 405102 582938 405134 583174
rect 404514 582854 405134 582938
rect 404514 582618 404546 582854
rect 404782 582618 404866 582854
rect 405102 582618 405134 582854
rect 404514 547174 405134 582618
rect 404514 546938 404546 547174
rect 404782 546938 404866 547174
rect 405102 546938 405134 547174
rect 404514 546854 405134 546938
rect 404514 546618 404546 546854
rect 404782 546618 404866 546854
rect 405102 546618 405134 546854
rect 404514 511174 405134 546618
rect 404514 510938 404546 511174
rect 404782 510938 404866 511174
rect 405102 510938 405134 511174
rect 404514 510854 405134 510938
rect 404514 510618 404546 510854
rect 404782 510618 404866 510854
rect 405102 510618 405134 510854
rect 404514 475174 405134 510618
rect 404514 474938 404546 475174
rect 404782 474938 404866 475174
rect 405102 474938 405134 475174
rect 404514 474854 405134 474938
rect 404514 474618 404546 474854
rect 404782 474618 404866 474854
rect 405102 474618 405134 474854
rect 404514 439174 405134 474618
rect 404514 438938 404546 439174
rect 404782 438938 404866 439174
rect 405102 438938 405134 439174
rect 404514 438854 405134 438938
rect 404514 438618 404546 438854
rect 404782 438618 404866 438854
rect 405102 438618 405134 438854
rect 404514 403174 405134 438618
rect 404514 402938 404546 403174
rect 404782 402938 404866 403174
rect 405102 402938 405134 403174
rect 404514 402854 405134 402938
rect 404514 402618 404546 402854
rect 404782 402618 404866 402854
rect 405102 402618 405134 402854
rect 404514 367174 405134 402618
rect 404514 366938 404546 367174
rect 404782 366938 404866 367174
rect 405102 366938 405134 367174
rect 404514 366854 405134 366938
rect 404514 366618 404546 366854
rect 404782 366618 404866 366854
rect 405102 366618 405134 366854
rect 404514 331174 405134 366618
rect 404514 330938 404546 331174
rect 404782 330938 404866 331174
rect 405102 330938 405134 331174
rect 404514 330854 405134 330938
rect 404514 330618 404546 330854
rect 404782 330618 404866 330854
rect 405102 330618 405134 330854
rect 404514 295174 405134 330618
rect 404514 294938 404546 295174
rect 404782 294938 404866 295174
rect 405102 294938 405134 295174
rect 404514 294854 405134 294938
rect 404514 294618 404546 294854
rect 404782 294618 404866 294854
rect 405102 294618 405134 294854
rect 404514 259174 405134 294618
rect 404514 258938 404546 259174
rect 404782 258938 404866 259174
rect 405102 258938 405134 259174
rect 404514 258854 405134 258938
rect 404514 258618 404546 258854
rect 404782 258618 404866 258854
rect 405102 258618 405134 258854
rect 404514 223174 405134 258618
rect 404514 222938 404546 223174
rect 404782 222938 404866 223174
rect 405102 222938 405134 223174
rect 404514 222854 405134 222938
rect 404514 222618 404546 222854
rect 404782 222618 404866 222854
rect 405102 222618 405134 222854
rect 404514 187174 405134 222618
rect 404514 186938 404546 187174
rect 404782 186938 404866 187174
rect 405102 186938 405134 187174
rect 404514 186854 405134 186938
rect 404514 186618 404546 186854
rect 404782 186618 404866 186854
rect 405102 186618 405134 186854
rect 404514 151174 405134 186618
rect 404514 150938 404546 151174
rect 404782 150938 404866 151174
rect 405102 150938 405134 151174
rect 404514 150854 405134 150938
rect 404514 150618 404546 150854
rect 404782 150618 404866 150854
rect 405102 150618 405134 150854
rect 404514 115174 405134 150618
rect 404514 114938 404546 115174
rect 404782 114938 404866 115174
rect 405102 114938 405134 115174
rect 404514 114854 405134 114938
rect 404514 114618 404546 114854
rect 404782 114618 404866 114854
rect 405102 114618 405134 114854
rect 404514 79174 405134 114618
rect 404514 78938 404546 79174
rect 404782 78938 404866 79174
rect 405102 78938 405134 79174
rect 404514 78854 405134 78938
rect 404514 78618 404546 78854
rect 404782 78618 404866 78854
rect 405102 78618 405134 78854
rect 404514 43174 405134 78618
rect 404514 42938 404546 43174
rect 404782 42938 404866 43174
rect 405102 42938 405134 43174
rect 404514 42854 405134 42938
rect 404514 42618 404546 42854
rect 404782 42618 404866 42854
rect 405102 42618 405134 42854
rect 404514 7174 405134 42618
rect 404514 6938 404546 7174
rect 404782 6938 404866 7174
rect 405102 6938 405134 7174
rect 404514 6854 405134 6938
rect 404514 6618 404546 6854
rect 404782 6618 404866 6854
rect 405102 6618 405134 6854
rect 404514 -2266 405134 6618
rect 404514 -2502 404546 -2266
rect 404782 -2502 404866 -2266
rect 405102 -2502 405134 -2266
rect 404514 -2586 405134 -2502
rect 404514 -2822 404546 -2586
rect 404782 -2822 404866 -2586
rect 405102 -2822 405134 -2586
rect 404514 -3814 405134 -2822
rect 408234 694894 408854 708122
rect 408234 694658 408266 694894
rect 408502 694658 408586 694894
rect 408822 694658 408854 694894
rect 408234 694574 408854 694658
rect 408234 694338 408266 694574
rect 408502 694338 408586 694574
rect 408822 694338 408854 694574
rect 408234 658894 408854 694338
rect 408234 658658 408266 658894
rect 408502 658658 408586 658894
rect 408822 658658 408854 658894
rect 408234 658574 408854 658658
rect 408234 658338 408266 658574
rect 408502 658338 408586 658574
rect 408822 658338 408854 658574
rect 408234 622894 408854 658338
rect 408234 622658 408266 622894
rect 408502 622658 408586 622894
rect 408822 622658 408854 622894
rect 408234 622574 408854 622658
rect 408234 622338 408266 622574
rect 408502 622338 408586 622574
rect 408822 622338 408854 622574
rect 408234 586894 408854 622338
rect 408234 586658 408266 586894
rect 408502 586658 408586 586894
rect 408822 586658 408854 586894
rect 408234 586574 408854 586658
rect 408234 586338 408266 586574
rect 408502 586338 408586 586574
rect 408822 586338 408854 586574
rect 408234 550894 408854 586338
rect 408234 550658 408266 550894
rect 408502 550658 408586 550894
rect 408822 550658 408854 550894
rect 408234 550574 408854 550658
rect 408234 550338 408266 550574
rect 408502 550338 408586 550574
rect 408822 550338 408854 550574
rect 408234 514894 408854 550338
rect 408234 514658 408266 514894
rect 408502 514658 408586 514894
rect 408822 514658 408854 514894
rect 408234 514574 408854 514658
rect 408234 514338 408266 514574
rect 408502 514338 408586 514574
rect 408822 514338 408854 514574
rect 408234 478894 408854 514338
rect 408234 478658 408266 478894
rect 408502 478658 408586 478894
rect 408822 478658 408854 478894
rect 408234 478574 408854 478658
rect 408234 478338 408266 478574
rect 408502 478338 408586 478574
rect 408822 478338 408854 478574
rect 408234 442894 408854 478338
rect 408234 442658 408266 442894
rect 408502 442658 408586 442894
rect 408822 442658 408854 442894
rect 408234 442574 408854 442658
rect 408234 442338 408266 442574
rect 408502 442338 408586 442574
rect 408822 442338 408854 442574
rect 408234 406894 408854 442338
rect 408234 406658 408266 406894
rect 408502 406658 408586 406894
rect 408822 406658 408854 406894
rect 408234 406574 408854 406658
rect 408234 406338 408266 406574
rect 408502 406338 408586 406574
rect 408822 406338 408854 406574
rect 408234 370894 408854 406338
rect 408234 370658 408266 370894
rect 408502 370658 408586 370894
rect 408822 370658 408854 370894
rect 408234 370574 408854 370658
rect 408234 370338 408266 370574
rect 408502 370338 408586 370574
rect 408822 370338 408854 370574
rect 408234 334894 408854 370338
rect 408234 334658 408266 334894
rect 408502 334658 408586 334894
rect 408822 334658 408854 334894
rect 408234 334574 408854 334658
rect 408234 334338 408266 334574
rect 408502 334338 408586 334574
rect 408822 334338 408854 334574
rect 408234 298894 408854 334338
rect 408234 298658 408266 298894
rect 408502 298658 408586 298894
rect 408822 298658 408854 298894
rect 408234 298574 408854 298658
rect 408234 298338 408266 298574
rect 408502 298338 408586 298574
rect 408822 298338 408854 298574
rect 408234 262894 408854 298338
rect 408234 262658 408266 262894
rect 408502 262658 408586 262894
rect 408822 262658 408854 262894
rect 408234 262574 408854 262658
rect 408234 262338 408266 262574
rect 408502 262338 408586 262574
rect 408822 262338 408854 262574
rect 408234 226894 408854 262338
rect 408234 226658 408266 226894
rect 408502 226658 408586 226894
rect 408822 226658 408854 226894
rect 408234 226574 408854 226658
rect 408234 226338 408266 226574
rect 408502 226338 408586 226574
rect 408822 226338 408854 226574
rect 408234 190894 408854 226338
rect 408234 190658 408266 190894
rect 408502 190658 408586 190894
rect 408822 190658 408854 190894
rect 408234 190574 408854 190658
rect 408234 190338 408266 190574
rect 408502 190338 408586 190574
rect 408822 190338 408854 190574
rect 408234 154894 408854 190338
rect 408234 154658 408266 154894
rect 408502 154658 408586 154894
rect 408822 154658 408854 154894
rect 408234 154574 408854 154658
rect 408234 154338 408266 154574
rect 408502 154338 408586 154574
rect 408822 154338 408854 154574
rect 408234 118894 408854 154338
rect 408234 118658 408266 118894
rect 408502 118658 408586 118894
rect 408822 118658 408854 118894
rect 408234 118574 408854 118658
rect 408234 118338 408266 118574
rect 408502 118338 408586 118574
rect 408822 118338 408854 118574
rect 408234 82894 408854 118338
rect 408234 82658 408266 82894
rect 408502 82658 408586 82894
rect 408822 82658 408854 82894
rect 408234 82574 408854 82658
rect 408234 82338 408266 82574
rect 408502 82338 408586 82574
rect 408822 82338 408854 82574
rect 408234 46894 408854 82338
rect 408234 46658 408266 46894
rect 408502 46658 408586 46894
rect 408822 46658 408854 46894
rect 408234 46574 408854 46658
rect 408234 46338 408266 46574
rect 408502 46338 408586 46574
rect 408822 46338 408854 46574
rect 408234 10894 408854 46338
rect 408234 10658 408266 10894
rect 408502 10658 408586 10894
rect 408822 10658 408854 10894
rect 408234 10574 408854 10658
rect 408234 10338 408266 10574
rect 408502 10338 408586 10574
rect 408822 10338 408854 10574
rect 408234 -4186 408854 10338
rect 410794 705798 411414 705830
rect 410794 705562 410826 705798
rect 411062 705562 411146 705798
rect 411382 705562 411414 705798
rect 410794 705478 411414 705562
rect 410794 705242 410826 705478
rect 411062 705242 411146 705478
rect 411382 705242 411414 705478
rect 410794 669454 411414 705242
rect 410794 669218 410826 669454
rect 411062 669218 411146 669454
rect 411382 669218 411414 669454
rect 410794 669134 411414 669218
rect 410794 668898 410826 669134
rect 411062 668898 411146 669134
rect 411382 668898 411414 669134
rect 410794 633454 411414 668898
rect 410794 633218 410826 633454
rect 411062 633218 411146 633454
rect 411382 633218 411414 633454
rect 410794 633134 411414 633218
rect 410794 632898 410826 633134
rect 411062 632898 411146 633134
rect 411382 632898 411414 633134
rect 410794 597454 411414 632898
rect 410794 597218 410826 597454
rect 411062 597218 411146 597454
rect 411382 597218 411414 597454
rect 410794 597134 411414 597218
rect 410794 596898 410826 597134
rect 411062 596898 411146 597134
rect 411382 596898 411414 597134
rect 410794 561454 411414 596898
rect 410794 561218 410826 561454
rect 411062 561218 411146 561454
rect 411382 561218 411414 561454
rect 410794 561134 411414 561218
rect 410794 560898 410826 561134
rect 411062 560898 411146 561134
rect 411382 560898 411414 561134
rect 410794 525454 411414 560898
rect 410794 525218 410826 525454
rect 411062 525218 411146 525454
rect 411382 525218 411414 525454
rect 410794 525134 411414 525218
rect 410794 524898 410826 525134
rect 411062 524898 411146 525134
rect 411382 524898 411414 525134
rect 410794 489454 411414 524898
rect 410794 489218 410826 489454
rect 411062 489218 411146 489454
rect 411382 489218 411414 489454
rect 410794 489134 411414 489218
rect 410794 488898 410826 489134
rect 411062 488898 411146 489134
rect 411382 488898 411414 489134
rect 410794 453454 411414 488898
rect 410794 453218 410826 453454
rect 411062 453218 411146 453454
rect 411382 453218 411414 453454
rect 410794 453134 411414 453218
rect 410794 452898 410826 453134
rect 411062 452898 411146 453134
rect 411382 452898 411414 453134
rect 410794 417454 411414 452898
rect 410794 417218 410826 417454
rect 411062 417218 411146 417454
rect 411382 417218 411414 417454
rect 410794 417134 411414 417218
rect 410794 416898 410826 417134
rect 411062 416898 411146 417134
rect 411382 416898 411414 417134
rect 410794 381454 411414 416898
rect 410794 381218 410826 381454
rect 411062 381218 411146 381454
rect 411382 381218 411414 381454
rect 410794 381134 411414 381218
rect 410794 380898 410826 381134
rect 411062 380898 411146 381134
rect 411382 380898 411414 381134
rect 410794 345454 411414 380898
rect 410794 345218 410826 345454
rect 411062 345218 411146 345454
rect 411382 345218 411414 345454
rect 410794 345134 411414 345218
rect 410794 344898 410826 345134
rect 411062 344898 411146 345134
rect 411382 344898 411414 345134
rect 410794 309454 411414 344898
rect 410794 309218 410826 309454
rect 411062 309218 411146 309454
rect 411382 309218 411414 309454
rect 410794 309134 411414 309218
rect 410794 308898 410826 309134
rect 411062 308898 411146 309134
rect 411382 308898 411414 309134
rect 410794 273454 411414 308898
rect 410794 273218 410826 273454
rect 411062 273218 411146 273454
rect 411382 273218 411414 273454
rect 410794 273134 411414 273218
rect 410794 272898 410826 273134
rect 411062 272898 411146 273134
rect 411382 272898 411414 273134
rect 410794 237454 411414 272898
rect 410794 237218 410826 237454
rect 411062 237218 411146 237454
rect 411382 237218 411414 237454
rect 410794 237134 411414 237218
rect 410794 236898 410826 237134
rect 411062 236898 411146 237134
rect 411382 236898 411414 237134
rect 410794 201454 411414 236898
rect 410794 201218 410826 201454
rect 411062 201218 411146 201454
rect 411382 201218 411414 201454
rect 410794 201134 411414 201218
rect 410794 200898 410826 201134
rect 411062 200898 411146 201134
rect 411382 200898 411414 201134
rect 410794 165454 411414 200898
rect 410794 165218 410826 165454
rect 411062 165218 411146 165454
rect 411382 165218 411414 165454
rect 410794 165134 411414 165218
rect 410794 164898 410826 165134
rect 411062 164898 411146 165134
rect 411382 164898 411414 165134
rect 410794 129454 411414 164898
rect 410794 129218 410826 129454
rect 411062 129218 411146 129454
rect 411382 129218 411414 129454
rect 410794 129134 411414 129218
rect 410794 128898 410826 129134
rect 411062 128898 411146 129134
rect 411382 128898 411414 129134
rect 410794 93454 411414 128898
rect 410794 93218 410826 93454
rect 411062 93218 411146 93454
rect 411382 93218 411414 93454
rect 410794 93134 411414 93218
rect 410794 92898 410826 93134
rect 411062 92898 411146 93134
rect 411382 92898 411414 93134
rect 410794 57454 411414 92898
rect 410794 57218 410826 57454
rect 411062 57218 411146 57454
rect 411382 57218 411414 57454
rect 410794 57134 411414 57218
rect 410794 56898 410826 57134
rect 411062 56898 411146 57134
rect 411382 56898 411414 57134
rect 410794 21454 411414 56898
rect 410794 21218 410826 21454
rect 411062 21218 411146 21454
rect 411382 21218 411414 21454
rect 410794 21134 411414 21218
rect 410794 20898 410826 21134
rect 411062 20898 411146 21134
rect 411382 20898 411414 21134
rect 410794 -1306 411414 20898
rect 410794 -1542 410826 -1306
rect 411062 -1542 411146 -1306
rect 411382 -1542 411414 -1306
rect 410794 -1626 411414 -1542
rect 410794 -1862 410826 -1626
rect 411062 -1862 411146 -1626
rect 411382 -1862 411414 -1626
rect 410794 -1894 411414 -1862
rect 411954 698614 412574 710042
rect 421954 711558 422574 711590
rect 421954 711322 421986 711558
rect 422222 711322 422306 711558
rect 422542 711322 422574 711558
rect 421954 711238 422574 711322
rect 421954 711002 421986 711238
rect 422222 711002 422306 711238
rect 422542 711002 422574 711238
rect 418234 709638 418854 709670
rect 418234 709402 418266 709638
rect 418502 709402 418586 709638
rect 418822 709402 418854 709638
rect 418234 709318 418854 709402
rect 418234 709082 418266 709318
rect 418502 709082 418586 709318
rect 418822 709082 418854 709318
rect 411954 698378 411986 698614
rect 412222 698378 412306 698614
rect 412542 698378 412574 698614
rect 411954 698294 412574 698378
rect 411954 698058 411986 698294
rect 412222 698058 412306 698294
rect 412542 698058 412574 698294
rect 411954 662614 412574 698058
rect 411954 662378 411986 662614
rect 412222 662378 412306 662614
rect 412542 662378 412574 662614
rect 411954 662294 412574 662378
rect 411954 662058 411986 662294
rect 412222 662058 412306 662294
rect 412542 662058 412574 662294
rect 411954 626614 412574 662058
rect 411954 626378 411986 626614
rect 412222 626378 412306 626614
rect 412542 626378 412574 626614
rect 411954 626294 412574 626378
rect 411954 626058 411986 626294
rect 412222 626058 412306 626294
rect 412542 626058 412574 626294
rect 411954 590614 412574 626058
rect 411954 590378 411986 590614
rect 412222 590378 412306 590614
rect 412542 590378 412574 590614
rect 411954 590294 412574 590378
rect 411954 590058 411986 590294
rect 412222 590058 412306 590294
rect 412542 590058 412574 590294
rect 411954 554614 412574 590058
rect 411954 554378 411986 554614
rect 412222 554378 412306 554614
rect 412542 554378 412574 554614
rect 411954 554294 412574 554378
rect 411954 554058 411986 554294
rect 412222 554058 412306 554294
rect 412542 554058 412574 554294
rect 411954 518614 412574 554058
rect 411954 518378 411986 518614
rect 412222 518378 412306 518614
rect 412542 518378 412574 518614
rect 411954 518294 412574 518378
rect 411954 518058 411986 518294
rect 412222 518058 412306 518294
rect 412542 518058 412574 518294
rect 411954 482614 412574 518058
rect 411954 482378 411986 482614
rect 412222 482378 412306 482614
rect 412542 482378 412574 482614
rect 411954 482294 412574 482378
rect 411954 482058 411986 482294
rect 412222 482058 412306 482294
rect 412542 482058 412574 482294
rect 411954 446614 412574 482058
rect 411954 446378 411986 446614
rect 412222 446378 412306 446614
rect 412542 446378 412574 446614
rect 411954 446294 412574 446378
rect 411954 446058 411986 446294
rect 412222 446058 412306 446294
rect 412542 446058 412574 446294
rect 411954 410614 412574 446058
rect 411954 410378 411986 410614
rect 412222 410378 412306 410614
rect 412542 410378 412574 410614
rect 411954 410294 412574 410378
rect 411954 410058 411986 410294
rect 412222 410058 412306 410294
rect 412542 410058 412574 410294
rect 411954 374614 412574 410058
rect 411954 374378 411986 374614
rect 412222 374378 412306 374614
rect 412542 374378 412574 374614
rect 411954 374294 412574 374378
rect 411954 374058 411986 374294
rect 412222 374058 412306 374294
rect 412542 374058 412574 374294
rect 411954 338614 412574 374058
rect 411954 338378 411986 338614
rect 412222 338378 412306 338614
rect 412542 338378 412574 338614
rect 411954 338294 412574 338378
rect 411954 338058 411986 338294
rect 412222 338058 412306 338294
rect 412542 338058 412574 338294
rect 411954 302614 412574 338058
rect 411954 302378 411986 302614
rect 412222 302378 412306 302614
rect 412542 302378 412574 302614
rect 411954 302294 412574 302378
rect 411954 302058 411986 302294
rect 412222 302058 412306 302294
rect 412542 302058 412574 302294
rect 411954 266614 412574 302058
rect 411954 266378 411986 266614
rect 412222 266378 412306 266614
rect 412542 266378 412574 266614
rect 411954 266294 412574 266378
rect 411954 266058 411986 266294
rect 412222 266058 412306 266294
rect 412542 266058 412574 266294
rect 411954 230614 412574 266058
rect 411954 230378 411986 230614
rect 412222 230378 412306 230614
rect 412542 230378 412574 230614
rect 411954 230294 412574 230378
rect 411954 230058 411986 230294
rect 412222 230058 412306 230294
rect 412542 230058 412574 230294
rect 411954 194614 412574 230058
rect 411954 194378 411986 194614
rect 412222 194378 412306 194614
rect 412542 194378 412574 194614
rect 411954 194294 412574 194378
rect 411954 194058 411986 194294
rect 412222 194058 412306 194294
rect 412542 194058 412574 194294
rect 411954 158614 412574 194058
rect 411954 158378 411986 158614
rect 412222 158378 412306 158614
rect 412542 158378 412574 158614
rect 411954 158294 412574 158378
rect 411954 158058 411986 158294
rect 412222 158058 412306 158294
rect 412542 158058 412574 158294
rect 411954 122614 412574 158058
rect 411954 122378 411986 122614
rect 412222 122378 412306 122614
rect 412542 122378 412574 122614
rect 411954 122294 412574 122378
rect 411954 122058 411986 122294
rect 412222 122058 412306 122294
rect 412542 122058 412574 122294
rect 411954 86614 412574 122058
rect 411954 86378 411986 86614
rect 412222 86378 412306 86614
rect 412542 86378 412574 86614
rect 411954 86294 412574 86378
rect 411954 86058 411986 86294
rect 412222 86058 412306 86294
rect 412542 86058 412574 86294
rect 411954 50614 412574 86058
rect 411954 50378 411986 50614
rect 412222 50378 412306 50614
rect 412542 50378 412574 50614
rect 411954 50294 412574 50378
rect 411954 50058 411986 50294
rect 412222 50058 412306 50294
rect 412542 50058 412574 50294
rect 411954 14614 412574 50058
rect 411954 14378 411986 14614
rect 412222 14378 412306 14614
rect 412542 14378 412574 14614
rect 411954 14294 412574 14378
rect 411954 14058 411986 14294
rect 412222 14058 412306 14294
rect 412542 14058 412574 14294
rect 408234 -4422 408266 -4186
rect 408502 -4422 408586 -4186
rect 408822 -4422 408854 -4186
rect 408234 -4506 408854 -4422
rect 408234 -4742 408266 -4506
rect 408502 -4742 408586 -4506
rect 408822 -4742 408854 -4506
rect 408234 -5734 408854 -4742
rect 401954 -7302 401986 -7066
rect 402222 -7302 402306 -7066
rect 402542 -7302 402574 -7066
rect 401954 -7386 402574 -7302
rect 401954 -7622 401986 -7386
rect 402222 -7622 402306 -7386
rect 402542 -7622 402574 -7386
rect 401954 -7654 402574 -7622
rect 411954 -6106 412574 14058
rect 414514 707718 415134 707750
rect 414514 707482 414546 707718
rect 414782 707482 414866 707718
rect 415102 707482 415134 707718
rect 414514 707398 415134 707482
rect 414514 707162 414546 707398
rect 414782 707162 414866 707398
rect 415102 707162 415134 707398
rect 414514 673174 415134 707162
rect 414514 672938 414546 673174
rect 414782 672938 414866 673174
rect 415102 672938 415134 673174
rect 414514 672854 415134 672938
rect 414514 672618 414546 672854
rect 414782 672618 414866 672854
rect 415102 672618 415134 672854
rect 414514 637174 415134 672618
rect 414514 636938 414546 637174
rect 414782 636938 414866 637174
rect 415102 636938 415134 637174
rect 414514 636854 415134 636938
rect 414514 636618 414546 636854
rect 414782 636618 414866 636854
rect 415102 636618 415134 636854
rect 414514 601174 415134 636618
rect 414514 600938 414546 601174
rect 414782 600938 414866 601174
rect 415102 600938 415134 601174
rect 414514 600854 415134 600938
rect 414514 600618 414546 600854
rect 414782 600618 414866 600854
rect 415102 600618 415134 600854
rect 414514 565174 415134 600618
rect 414514 564938 414546 565174
rect 414782 564938 414866 565174
rect 415102 564938 415134 565174
rect 414514 564854 415134 564938
rect 414514 564618 414546 564854
rect 414782 564618 414866 564854
rect 415102 564618 415134 564854
rect 414514 529174 415134 564618
rect 414514 528938 414546 529174
rect 414782 528938 414866 529174
rect 415102 528938 415134 529174
rect 414514 528854 415134 528938
rect 414514 528618 414546 528854
rect 414782 528618 414866 528854
rect 415102 528618 415134 528854
rect 414514 493174 415134 528618
rect 414514 492938 414546 493174
rect 414782 492938 414866 493174
rect 415102 492938 415134 493174
rect 414514 492854 415134 492938
rect 414514 492618 414546 492854
rect 414782 492618 414866 492854
rect 415102 492618 415134 492854
rect 414514 457174 415134 492618
rect 414514 456938 414546 457174
rect 414782 456938 414866 457174
rect 415102 456938 415134 457174
rect 414514 456854 415134 456938
rect 414514 456618 414546 456854
rect 414782 456618 414866 456854
rect 415102 456618 415134 456854
rect 414514 421174 415134 456618
rect 414514 420938 414546 421174
rect 414782 420938 414866 421174
rect 415102 420938 415134 421174
rect 414514 420854 415134 420938
rect 414514 420618 414546 420854
rect 414782 420618 414866 420854
rect 415102 420618 415134 420854
rect 414514 385174 415134 420618
rect 414514 384938 414546 385174
rect 414782 384938 414866 385174
rect 415102 384938 415134 385174
rect 414514 384854 415134 384938
rect 414514 384618 414546 384854
rect 414782 384618 414866 384854
rect 415102 384618 415134 384854
rect 414514 349174 415134 384618
rect 414514 348938 414546 349174
rect 414782 348938 414866 349174
rect 415102 348938 415134 349174
rect 414514 348854 415134 348938
rect 414514 348618 414546 348854
rect 414782 348618 414866 348854
rect 415102 348618 415134 348854
rect 414514 313174 415134 348618
rect 414514 312938 414546 313174
rect 414782 312938 414866 313174
rect 415102 312938 415134 313174
rect 414514 312854 415134 312938
rect 414514 312618 414546 312854
rect 414782 312618 414866 312854
rect 415102 312618 415134 312854
rect 414514 277174 415134 312618
rect 414514 276938 414546 277174
rect 414782 276938 414866 277174
rect 415102 276938 415134 277174
rect 414514 276854 415134 276938
rect 414514 276618 414546 276854
rect 414782 276618 414866 276854
rect 415102 276618 415134 276854
rect 414514 241174 415134 276618
rect 414514 240938 414546 241174
rect 414782 240938 414866 241174
rect 415102 240938 415134 241174
rect 414514 240854 415134 240938
rect 414514 240618 414546 240854
rect 414782 240618 414866 240854
rect 415102 240618 415134 240854
rect 414514 205174 415134 240618
rect 414514 204938 414546 205174
rect 414782 204938 414866 205174
rect 415102 204938 415134 205174
rect 414514 204854 415134 204938
rect 414514 204618 414546 204854
rect 414782 204618 414866 204854
rect 415102 204618 415134 204854
rect 414514 169174 415134 204618
rect 414514 168938 414546 169174
rect 414782 168938 414866 169174
rect 415102 168938 415134 169174
rect 414514 168854 415134 168938
rect 414514 168618 414546 168854
rect 414782 168618 414866 168854
rect 415102 168618 415134 168854
rect 414514 133174 415134 168618
rect 414514 132938 414546 133174
rect 414782 132938 414866 133174
rect 415102 132938 415134 133174
rect 414514 132854 415134 132938
rect 414514 132618 414546 132854
rect 414782 132618 414866 132854
rect 415102 132618 415134 132854
rect 414514 97174 415134 132618
rect 414514 96938 414546 97174
rect 414782 96938 414866 97174
rect 415102 96938 415134 97174
rect 414514 96854 415134 96938
rect 414514 96618 414546 96854
rect 414782 96618 414866 96854
rect 415102 96618 415134 96854
rect 414514 61174 415134 96618
rect 414514 60938 414546 61174
rect 414782 60938 414866 61174
rect 415102 60938 415134 61174
rect 414514 60854 415134 60938
rect 414514 60618 414546 60854
rect 414782 60618 414866 60854
rect 415102 60618 415134 60854
rect 414514 25174 415134 60618
rect 414514 24938 414546 25174
rect 414782 24938 414866 25174
rect 415102 24938 415134 25174
rect 414514 24854 415134 24938
rect 414514 24618 414546 24854
rect 414782 24618 414866 24854
rect 415102 24618 415134 24854
rect 414514 -3226 415134 24618
rect 414514 -3462 414546 -3226
rect 414782 -3462 414866 -3226
rect 415102 -3462 415134 -3226
rect 414514 -3546 415134 -3462
rect 414514 -3782 414546 -3546
rect 414782 -3782 414866 -3546
rect 415102 -3782 415134 -3546
rect 414514 -3814 415134 -3782
rect 418234 676894 418854 709082
rect 418234 676658 418266 676894
rect 418502 676658 418586 676894
rect 418822 676658 418854 676894
rect 418234 676574 418854 676658
rect 418234 676338 418266 676574
rect 418502 676338 418586 676574
rect 418822 676338 418854 676574
rect 418234 640894 418854 676338
rect 418234 640658 418266 640894
rect 418502 640658 418586 640894
rect 418822 640658 418854 640894
rect 418234 640574 418854 640658
rect 418234 640338 418266 640574
rect 418502 640338 418586 640574
rect 418822 640338 418854 640574
rect 418234 604894 418854 640338
rect 418234 604658 418266 604894
rect 418502 604658 418586 604894
rect 418822 604658 418854 604894
rect 418234 604574 418854 604658
rect 418234 604338 418266 604574
rect 418502 604338 418586 604574
rect 418822 604338 418854 604574
rect 418234 568894 418854 604338
rect 418234 568658 418266 568894
rect 418502 568658 418586 568894
rect 418822 568658 418854 568894
rect 418234 568574 418854 568658
rect 418234 568338 418266 568574
rect 418502 568338 418586 568574
rect 418822 568338 418854 568574
rect 418234 532894 418854 568338
rect 418234 532658 418266 532894
rect 418502 532658 418586 532894
rect 418822 532658 418854 532894
rect 418234 532574 418854 532658
rect 418234 532338 418266 532574
rect 418502 532338 418586 532574
rect 418822 532338 418854 532574
rect 418234 496894 418854 532338
rect 418234 496658 418266 496894
rect 418502 496658 418586 496894
rect 418822 496658 418854 496894
rect 418234 496574 418854 496658
rect 418234 496338 418266 496574
rect 418502 496338 418586 496574
rect 418822 496338 418854 496574
rect 418234 460894 418854 496338
rect 418234 460658 418266 460894
rect 418502 460658 418586 460894
rect 418822 460658 418854 460894
rect 418234 460574 418854 460658
rect 418234 460338 418266 460574
rect 418502 460338 418586 460574
rect 418822 460338 418854 460574
rect 418234 424894 418854 460338
rect 418234 424658 418266 424894
rect 418502 424658 418586 424894
rect 418822 424658 418854 424894
rect 418234 424574 418854 424658
rect 418234 424338 418266 424574
rect 418502 424338 418586 424574
rect 418822 424338 418854 424574
rect 418234 388894 418854 424338
rect 418234 388658 418266 388894
rect 418502 388658 418586 388894
rect 418822 388658 418854 388894
rect 418234 388574 418854 388658
rect 418234 388338 418266 388574
rect 418502 388338 418586 388574
rect 418822 388338 418854 388574
rect 418234 352894 418854 388338
rect 418234 352658 418266 352894
rect 418502 352658 418586 352894
rect 418822 352658 418854 352894
rect 418234 352574 418854 352658
rect 418234 352338 418266 352574
rect 418502 352338 418586 352574
rect 418822 352338 418854 352574
rect 418234 316894 418854 352338
rect 418234 316658 418266 316894
rect 418502 316658 418586 316894
rect 418822 316658 418854 316894
rect 418234 316574 418854 316658
rect 418234 316338 418266 316574
rect 418502 316338 418586 316574
rect 418822 316338 418854 316574
rect 418234 280894 418854 316338
rect 418234 280658 418266 280894
rect 418502 280658 418586 280894
rect 418822 280658 418854 280894
rect 418234 280574 418854 280658
rect 418234 280338 418266 280574
rect 418502 280338 418586 280574
rect 418822 280338 418854 280574
rect 418234 244894 418854 280338
rect 418234 244658 418266 244894
rect 418502 244658 418586 244894
rect 418822 244658 418854 244894
rect 418234 244574 418854 244658
rect 418234 244338 418266 244574
rect 418502 244338 418586 244574
rect 418822 244338 418854 244574
rect 418234 208894 418854 244338
rect 418234 208658 418266 208894
rect 418502 208658 418586 208894
rect 418822 208658 418854 208894
rect 418234 208574 418854 208658
rect 418234 208338 418266 208574
rect 418502 208338 418586 208574
rect 418822 208338 418854 208574
rect 418234 172894 418854 208338
rect 418234 172658 418266 172894
rect 418502 172658 418586 172894
rect 418822 172658 418854 172894
rect 418234 172574 418854 172658
rect 418234 172338 418266 172574
rect 418502 172338 418586 172574
rect 418822 172338 418854 172574
rect 418234 136894 418854 172338
rect 418234 136658 418266 136894
rect 418502 136658 418586 136894
rect 418822 136658 418854 136894
rect 418234 136574 418854 136658
rect 418234 136338 418266 136574
rect 418502 136338 418586 136574
rect 418822 136338 418854 136574
rect 418234 100894 418854 136338
rect 418234 100658 418266 100894
rect 418502 100658 418586 100894
rect 418822 100658 418854 100894
rect 418234 100574 418854 100658
rect 418234 100338 418266 100574
rect 418502 100338 418586 100574
rect 418822 100338 418854 100574
rect 418234 64894 418854 100338
rect 418234 64658 418266 64894
rect 418502 64658 418586 64894
rect 418822 64658 418854 64894
rect 418234 64574 418854 64658
rect 418234 64338 418266 64574
rect 418502 64338 418586 64574
rect 418822 64338 418854 64574
rect 418234 28894 418854 64338
rect 418234 28658 418266 28894
rect 418502 28658 418586 28894
rect 418822 28658 418854 28894
rect 418234 28574 418854 28658
rect 418234 28338 418266 28574
rect 418502 28338 418586 28574
rect 418822 28338 418854 28574
rect 418234 -5146 418854 28338
rect 420794 704838 421414 705830
rect 420794 704602 420826 704838
rect 421062 704602 421146 704838
rect 421382 704602 421414 704838
rect 420794 704518 421414 704602
rect 420794 704282 420826 704518
rect 421062 704282 421146 704518
rect 421382 704282 421414 704518
rect 420794 687454 421414 704282
rect 420794 687218 420826 687454
rect 421062 687218 421146 687454
rect 421382 687218 421414 687454
rect 420794 687134 421414 687218
rect 420794 686898 420826 687134
rect 421062 686898 421146 687134
rect 421382 686898 421414 687134
rect 420794 651454 421414 686898
rect 420794 651218 420826 651454
rect 421062 651218 421146 651454
rect 421382 651218 421414 651454
rect 420794 651134 421414 651218
rect 420794 650898 420826 651134
rect 421062 650898 421146 651134
rect 421382 650898 421414 651134
rect 420794 615454 421414 650898
rect 420794 615218 420826 615454
rect 421062 615218 421146 615454
rect 421382 615218 421414 615454
rect 420794 615134 421414 615218
rect 420794 614898 420826 615134
rect 421062 614898 421146 615134
rect 421382 614898 421414 615134
rect 420794 579454 421414 614898
rect 420794 579218 420826 579454
rect 421062 579218 421146 579454
rect 421382 579218 421414 579454
rect 420794 579134 421414 579218
rect 420794 578898 420826 579134
rect 421062 578898 421146 579134
rect 421382 578898 421414 579134
rect 420794 543454 421414 578898
rect 420794 543218 420826 543454
rect 421062 543218 421146 543454
rect 421382 543218 421414 543454
rect 420794 543134 421414 543218
rect 420794 542898 420826 543134
rect 421062 542898 421146 543134
rect 421382 542898 421414 543134
rect 420794 507454 421414 542898
rect 420794 507218 420826 507454
rect 421062 507218 421146 507454
rect 421382 507218 421414 507454
rect 420794 507134 421414 507218
rect 420794 506898 420826 507134
rect 421062 506898 421146 507134
rect 421382 506898 421414 507134
rect 420794 471454 421414 506898
rect 420794 471218 420826 471454
rect 421062 471218 421146 471454
rect 421382 471218 421414 471454
rect 420794 471134 421414 471218
rect 420794 470898 420826 471134
rect 421062 470898 421146 471134
rect 421382 470898 421414 471134
rect 420794 435454 421414 470898
rect 420794 435218 420826 435454
rect 421062 435218 421146 435454
rect 421382 435218 421414 435454
rect 420794 435134 421414 435218
rect 420794 434898 420826 435134
rect 421062 434898 421146 435134
rect 421382 434898 421414 435134
rect 420794 399454 421414 434898
rect 420794 399218 420826 399454
rect 421062 399218 421146 399454
rect 421382 399218 421414 399454
rect 420794 399134 421414 399218
rect 420794 398898 420826 399134
rect 421062 398898 421146 399134
rect 421382 398898 421414 399134
rect 420794 363454 421414 398898
rect 420794 363218 420826 363454
rect 421062 363218 421146 363454
rect 421382 363218 421414 363454
rect 420794 363134 421414 363218
rect 420794 362898 420826 363134
rect 421062 362898 421146 363134
rect 421382 362898 421414 363134
rect 420794 327454 421414 362898
rect 420794 327218 420826 327454
rect 421062 327218 421146 327454
rect 421382 327218 421414 327454
rect 420794 327134 421414 327218
rect 420794 326898 420826 327134
rect 421062 326898 421146 327134
rect 421382 326898 421414 327134
rect 420794 291454 421414 326898
rect 420794 291218 420826 291454
rect 421062 291218 421146 291454
rect 421382 291218 421414 291454
rect 420794 291134 421414 291218
rect 420794 290898 420826 291134
rect 421062 290898 421146 291134
rect 421382 290898 421414 291134
rect 420794 255454 421414 290898
rect 420794 255218 420826 255454
rect 421062 255218 421146 255454
rect 421382 255218 421414 255454
rect 420794 255134 421414 255218
rect 420794 254898 420826 255134
rect 421062 254898 421146 255134
rect 421382 254898 421414 255134
rect 420794 219454 421414 254898
rect 420794 219218 420826 219454
rect 421062 219218 421146 219454
rect 421382 219218 421414 219454
rect 420794 219134 421414 219218
rect 420794 218898 420826 219134
rect 421062 218898 421146 219134
rect 421382 218898 421414 219134
rect 420794 183454 421414 218898
rect 420794 183218 420826 183454
rect 421062 183218 421146 183454
rect 421382 183218 421414 183454
rect 420794 183134 421414 183218
rect 420794 182898 420826 183134
rect 421062 182898 421146 183134
rect 421382 182898 421414 183134
rect 420794 147454 421414 182898
rect 420794 147218 420826 147454
rect 421062 147218 421146 147454
rect 421382 147218 421414 147454
rect 420794 147134 421414 147218
rect 420794 146898 420826 147134
rect 421062 146898 421146 147134
rect 421382 146898 421414 147134
rect 420794 111454 421414 146898
rect 420794 111218 420826 111454
rect 421062 111218 421146 111454
rect 421382 111218 421414 111454
rect 420794 111134 421414 111218
rect 420794 110898 420826 111134
rect 421062 110898 421146 111134
rect 421382 110898 421414 111134
rect 420794 75454 421414 110898
rect 420794 75218 420826 75454
rect 421062 75218 421146 75454
rect 421382 75218 421414 75454
rect 420794 75134 421414 75218
rect 420794 74898 420826 75134
rect 421062 74898 421146 75134
rect 421382 74898 421414 75134
rect 420794 39454 421414 74898
rect 420794 39218 420826 39454
rect 421062 39218 421146 39454
rect 421382 39218 421414 39454
rect 420794 39134 421414 39218
rect 420794 38898 420826 39134
rect 421062 38898 421146 39134
rect 421382 38898 421414 39134
rect 420794 3454 421414 38898
rect 420794 3218 420826 3454
rect 421062 3218 421146 3454
rect 421382 3218 421414 3454
rect 420794 3134 421414 3218
rect 420794 2898 420826 3134
rect 421062 2898 421146 3134
rect 421382 2898 421414 3134
rect 420794 -346 421414 2898
rect 420794 -582 420826 -346
rect 421062 -582 421146 -346
rect 421382 -582 421414 -346
rect 420794 -666 421414 -582
rect 420794 -902 420826 -666
rect 421062 -902 421146 -666
rect 421382 -902 421414 -666
rect 420794 -1894 421414 -902
rect 421954 680614 422574 711002
rect 431954 710598 432574 711590
rect 431954 710362 431986 710598
rect 432222 710362 432306 710598
rect 432542 710362 432574 710598
rect 431954 710278 432574 710362
rect 431954 710042 431986 710278
rect 432222 710042 432306 710278
rect 432542 710042 432574 710278
rect 428234 708678 428854 709670
rect 428234 708442 428266 708678
rect 428502 708442 428586 708678
rect 428822 708442 428854 708678
rect 428234 708358 428854 708442
rect 428234 708122 428266 708358
rect 428502 708122 428586 708358
rect 428822 708122 428854 708358
rect 421954 680378 421986 680614
rect 422222 680378 422306 680614
rect 422542 680378 422574 680614
rect 421954 680294 422574 680378
rect 421954 680058 421986 680294
rect 422222 680058 422306 680294
rect 422542 680058 422574 680294
rect 421954 644614 422574 680058
rect 421954 644378 421986 644614
rect 422222 644378 422306 644614
rect 422542 644378 422574 644614
rect 421954 644294 422574 644378
rect 421954 644058 421986 644294
rect 422222 644058 422306 644294
rect 422542 644058 422574 644294
rect 421954 608614 422574 644058
rect 421954 608378 421986 608614
rect 422222 608378 422306 608614
rect 422542 608378 422574 608614
rect 421954 608294 422574 608378
rect 421954 608058 421986 608294
rect 422222 608058 422306 608294
rect 422542 608058 422574 608294
rect 421954 572614 422574 608058
rect 421954 572378 421986 572614
rect 422222 572378 422306 572614
rect 422542 572378 422574 572614
rect 421954 572294 422574 572378
rect 421954 572058 421986 572294
rect 422222 572058 422306 572294
rect 422542 572058 422574 572294
rect 421954 536614 422574 572058
rect 421954 536378 421986 536614
rect 422222 536378 422306 536614
rect 422542 536378 422574 536614
rect 421954 536294 422574 536378
rect 421954 536058 421986 536294
rect 422222 536058 422306 536294
rect 422542 536058 422574 536294
rect 421954 500614 422574 536058
rect 421954 500378 421986 500614
rect 422222 500378 422306 500614
rect 422542 500378 422574 500614
rect 421954 500294 422574 500378
rect 421954 500058 421986 500294
rect 422222 500058 422306 500294
rect 422542 500058 422574 500294
rect 421954 464614 422574 500058
rect 421954 464378 421986 464614
rect 422222 464378 422306 464614
rect 422542 464378 422574 464614
rect 421954 464294 422574 464378
rect 421954 464058 421986 464294
rect 422222 464058 422306 464294
rect 422542 464058 422574 464294
rect 421954 428614 422574 464058
rect 421954 428378 421986 428614
rect 422222 428378 422306 428614
rect 422542 428378 422574 428614
rect 421954 428294 422574 428378
rect 421954 428058 421986 428294
rect 422222 428058 422306 428294
rect 422542 428058 422574 428294
rect 421954 392614 422574 428058
rect 421954 392378 421986 392614
rect 422222 392378 422306 392614
rect 422542 392378 422574 392614
rect 421954 392294 422574 392378
rect 421954 392058 421986 392294
rect 422222 392058 422306 392294
rect 422542 392058 422574 392294
rect 421954 356614 422574 392058
rect 421954 356378 421986 356614
rect 422222 356378 422306 356614
rect 422542 356378 422574 356614
rect 421954 356294 422574 356378
rect 421954 356058 421986 356294
rect 422222 356058 422306 356294
rect 422542 356058 422574 356294
rect 421954 320614 422574 356058
rect 421954 320378 421986 320614
rect 422222 320378 422306 320614
rect 422542 320378 422574 320614
rect 421954 320294 422574 320378
rect 421954 320058 421986 320294
rect 422222 320058 422306 320294
rect 422542 320058 422574 320294
rect 421954 284614 422574 320058
rect 421954 284378 421986 284614
rect 422222 284378 422306 284614
rect 422542 284378 422574 284614
rect 421954 284294 422574 284378
rect 421954 284058 421986 284294
rect 422222 284058 422306 284294
rect 422542 284058 422574 284294
rect 421954 248614 422574 284058
rect 421954 248378 421986 248614
rect 422222 248378 422306 248614
rect 422542 248378 422574 248614
rect 421954 248294 422574 248378
rect 421954 248058 421986 248294
rect 422222 248058 422306 248294
rect 422542 248058 422574 248294
rect 421954 212614 422574 248058
rect 421954 212378 421986 212614
rect 422222 212378 422306 212614
rect 422542 212378 422574 212614
rect 421954 212294 422574 212378
rect 421954 212058 421986 212294
rect 422222 212058 422306 212294
rect 422542 212058 422574 212294
rect 421954 176614 422574 212058
rect 421954 176378 421986 176614
rect 422222 176378 422306 176614
rect 422542 176378 422574 176614
rect 421954 176294 422574 176378
rect 421954 176058 421986 176294
rect 422222 176058 422306 176294
rect 422542 176058 422574 176294
rect 421954 140614 422574 176058
rect 421954 140378 421986 140614
rect 422222 140378 422306 140614
rect 422542 140378 422574 140614
rect 421954 140294 422574 140378
rect 421954 140058 421986 140294
rect 422222 140058 422306 140294
rect 422542 140058 422574 140294
rect 421954 104614 422574 140058
rect 421954 104378 421986 104614
rect 422222 104378 422306 104614
rect 422542 104378 422574 104614
rect 421954 104294 422574 104378
rect 421954 104058 421986 104294
rect 422222 104058 422306 104294
rect 422542 104058 422574 104294
rect 421954 68614 422574 104058
rect 421954 68378 421986 68614
rect 422222 68378 422306 68614
rect 422542 68378 422574 68614
rect 421954 68294 422574 68378
rect 421954 68058 421986 68294
rect 422222 68058 422306 68294
rect 422542 68058 422574 68294
rect 421954 32614 422574 68058
rect 421954 32378 421986 32614
rect 422222 32378 422306 32614
rect 422542 32378 422574 32614
rect 421954 32294 422574 32378
rect 421954 32058 421986 32294
rect 422222 32058 422306 32294
rect 422542 32058 422574 32294
rect 418234 -5382 418266 -5146
rect 418502 -5382 418586 -5146
rect 418822 -5382 418854 -5146
rect 418234 -5466 418854 -5382
rect 418234 -5702 418266 -5466
rect 418502 -5702 418586 -5466
rect 418822 -5702 418854 -5466
rect 418234 -5734 418854 -5702
rect 411954 -6342 411986 -6106
rect 412222 -6342 412306 -6106
rect 412542 -6342 412574 -6106
rect 411954 -6426 412574 -6342
rect 411954 -6662 411986 -6426
rect 412222 -6662 412306 -6426
rect 412542 -6662 412574 -6426
rect 411954 -7654 412574 -6662
rect 421954 -7066 422574 32058
rect 424514 706758 425134 707750
rect 424514 706522 424546 706758
rect 424782 706522 424866 706758
rect 425102 706522 425134 706758
rect 424514 706438 425134 706522
rect 424514 706202 424546 706438
rect 424782 706202 424866 706438
rect 425102 706202 425134 706438
rect 424514 691174 425134 706202
rect 424514 690938 424546 691174
rect 424782 690938 424866 691174
rect 425102 690938 425134 691174
rect 424514 690854 425134 690938
rect 424514 690618 424546 690854
rect 424782 690618 424866 690854
rect 425102 690618 425134 690854
rect 424514 655174 425134 690618
rect 424514 654938 424546 655174
rect 424782 654938 424866 655174
rect 425102 654938 425134 655174
rect 424514 654854 425134 654938
rect 424514 654618 424546 654854
rect 424782 654618 424866 654854
rect 425102 654618 425134 654854
rect 424514 619174 425134 654618
rect 424514 618938 424546 619174
rect 424782 618938 424866 619174
rect 425102 618938 425134 619174
rect 424514 618854 425134 618938
rect 424514 618618 424546 618854
rect 424782 618618 424866 618854
rect 425102 618618 425134 618854
rect 424514 583174 425134 618618
rect 424514 582938 424546 583174
rect 424782 582938 424866 583174
rect 425102 582938 425134 583174
rect 424514 582854 425134 582938
rect 424514 582618 424546 582854
rect 424782 582618 424866 582854
rect 425102 582618 425134 582854
rect 424514 547174 425134 582618
rect 424514 546938 424546 547174
rect 424782 546938 424866 547174
rect 425102 546938 425134 547174
rect 424514 546854 425134 546938
rect 424514 546618 424546 546854
rect 424782 546618 424866 546854
rect 425102 546618 425134 546854
rect 424514 511174 425134 546618
rect 424514 510938 424546 511174
rect 424782 510938 424866 511174
rect 425102 510938 425134 511174
rect 424514 510854 425134 510938
rect 424514 510618 424546 510854
rect 424782 510618 424866 510854
rect 425102 510618 425134 510854
rect 424514 475174 425134 510618
rect 424514 474938 424546 475174
rect 424782 474938 424866 475174
rect 425102 474938 425134 475174
rect 424514 474854 425134 474938
rect 424514 474618 424546 474854
rect 424782 474618 424866 474854
rect 425102 474618 425134 474854
rect 424514 439174 425134 474618
rect 424514 438938 424546 439174
rect 424782 438938 424866 439174
rect 425102 438938 425134 439174
rect 424514 438854 425134 438938
rect 424514 438618 424546 438854
rect 424782 438618 424866 438854
rect 425102 438618 425134 438854
rect 424514 403174 425134 438618
rect 424514 402938 424546 403174
rect 424782 402938 424866 403174
rect 425102 402938 425134 403174
rect 424514 402854 425134 402938
rect 424514 402618 424546 402854
rect 424782 402618 424866 402854
rect 425102 402618 425134 402854
rect 424514 367174 425134 402618
rect 424514 366938 424546 367174
rect 424782 366938 424866 367174
rect 425102 366938 425134 367174
rect 424514 366854 425134 366938
rect 424514 366618 424546 366854
rect 424782 366618 424866 366854
rect 425102 366618 425134 366854
rect 424514 331174 425134 366618
rect 424514 330938 424546 331174
rect 424782 330938 424866 331174
rect 425102 330938 425134 331174
rect 424514 330854 425134 330938
rect 424514 330618 424546 330854
rect 424782 330618 424866 330854
rect 425102 330618 425134 330854
rect 424514 295174 425134 330618
rect 424514 294938 424546 295174
rect 424782 294938 424866 295174
rect 425102 294938 425134 295174
rect 424514 294854 425134 294938
rect 424514 294618 424546 294854
rect 424782 294618 424866 294854
rect 425102 294618 425134 294854
rect 424514 259174 425134 294618
rect 424514 258938 424546 259174
rect 424782 258938 424866 259174
rect 425102 258938 425134 259174
rect 424514 258854 425134 258938
rect 424514 258618 424546 258854
rect 424782 258618 424866 258854
rect 425102 258618 425134 258854
rect 424514 223174 425134 258618
rect 424514 222938 424546 223174
rect 424782 222938 424866 223174
rect 425102 222938 425134 223174
rect 424514 222854 425134 222938
rect 424514 222618 424546 222854
rect 424782 222618 424866 222854
rect 425102 222618 425134 222854
rect 424514 187174 425134 222618
rect 424514 186938 424546 187174
rect 424782 186938 424866 187174
rect 425102 186938 425134 187174
rect 424514 186854 425134 186938
rect 424514 186618 424546 186854
rect 424782 186618 424866 186854
rect 425102 186618 425134 186854
rect 424514 151174 425134 186618
rect 424514 150938 424546 151174
rect 424782 150938 424866 151174
rect 425102 150938 425134 151174
rect 424514 150854 425134 150938
rect 424514 150618 424546 150854
rect 424782 150618 424866 150854
rect 425102 150618 425134 150854
rect 424514 115174 425134 150618
rect 424514 114938 424546 115174
rect 424782 114938 424866 115174
rect 425102 114938 425134 115174
rect 424514 114854 425134 114938
rect 424514 114618 424546 114854
rect 424782 114618 424866 114854
rect 425102 114618 425134 114854
rect 424514 79174 425134 114618
rect 424514 78938 424546 79174
rect 424782 78938 424866 79174
rect 425102 78938 425134 79174
rect 424514 78854 425134 78938
rect 424514 78618 424546 78854
rect 424782 78618 424866 78854
rect 425102 78618 425134 78854
rect 424514 43174 425134 78618
rect 424514 42938 424546 43174
rect 424782 42938 424866 43174
rect 425102 42938 425134 43174
rect 424514 42854 425134 42938
rect 424514 42618 424546 42854
rect 424782 42618 424866 42854
rect 425102 42618 425134 42854
rect 424514 7174 425134 42618
rect 424514 6938 424546 7174
rect 424782 6938 424866 7174
rect 425102 6938 425134 7174
rect 424514 6854 425134 6938
rect 424514 6618 424546 6854
rect 424782 6618 424866 6854
rect 425102 6618 425134 6854
rect 424514 -2266 425134 6618
rect 424514 -2502 424546 -2266
rect 424782 -2502 424866 -2266
rect 425102 -2502 425134 -2266
rect 424514 -2586 425134 -2502
rect 424514 -2822 424546 -2586
rect 424782 -2822 424866 -2586
rect 425102 -2822 425134 -2586
rect 424514 -3814 425134 -2822
rect 428234 694894 428854 708122
rect 428234 694658 428266 694894
rect 428502 694658 428586 694894
rect 428822 694658 428854 694894
rect 428234 694574 428854 694658
rect 428234 694338 428266 694574
rect 428502 694338 428586 694574
rect 428822 694338 428854 694574
rect 428234 658894 428854 694338
rect 428234 658658 428266 658894
rect 428502 658658 428586 658894
rect 428822 658658 428854 658894
rect 428234 658574 428854 658658
rect 428234 658338 428266 658574
rect 428502 658338 428586 658574
rect 428822 658338 428854 658574
rect 428234 622894 428854 658338
rect 428234 622658 428266 622894
rect 428502 622658 428586 622894
rect 428822 622658 428854 622894
rect 428234 622574 428854 622658
rect 428234 622338 428266 622574
rect 428502 622338 428586 622574
rect 428822 622338 428854 622574
rect 428234 586894 428854 622338
rect 428234 586658 428266 586894
rect 428502 586658 428586 586894
rect 428822 586658 428854 586894
rect 428234 586574 428854 586658
rect 428234 586338 428266 586574
rect 428502 586338 428586 586574
rect 428822 586338 428854 586574
rect 428234 550894 428854 586338
rect 428234 550658 428266 550894
rect 428502 550658 428586 550894
rect 428822 550658 428854 550894
rect 428234 550574 428854 550658
rect 428234 550338 428266 550574
rect 428502 550338 428586 550574
rect 428822 550338 428854 550574
rect 428234 514894 428854 550338
rect 428234 514658 428266 514894
rect 428502 514658 428586 514894
rect 428822 514658 428854 514894
rect 428234 514574 428854 514658
rect 428234 514338 428266 514574
rect 428502 514338 428586 514574
rect 428822 514338 428854 514574
rect 428234 478894 428854 514338
rect 428234 478658 428266 478894
rect 428502 478658 428586 478894
rect 428822 478658 428854 478894
rect 428234 478574 428854 478658
rect 428234 478338 428266 478574
rect 428502 478338 428586 478574
rect 428822 478338 428854 478574
rect 428234 442894 428854 478338
rect 428234 442658 428266 442894
rect 428502 442658 428586 442894
rect 428822 442658 428854 442894
rect 428234 442574 428854 442658
rect 428234 442338 428266 442574
rect 428502 442338 428586 442574
rect 428822 442338 428854 442574
rect 428234 406894 428854 442338
rect 428234 406658 428266 406894
rect 428502 406658 428586 406894
rect 428822 406658 428854 406894
rect 428234 406574 428854 406658
rect 428234 406338 428266 406574
rect 428502 406338 428586 406574
rect 428822 406338 428854 406574
rect 428234 370894 428854 406338
rect 428234 370658 428266 370894
rect 428502 370658 428586 370894
rect 428822 370658 428854 370894
rect 428234 370574 428854 370658
rect 428234 370338 428266 370574
rect 428502 370338 428586 370574
rect 428822 370338 428854 370574
rect 428234 334894 428854 370338
rect 428234 334658 428266 334894
rect 428502 334658 428586 334894
rect 428822 334658 428854 334894
rect 428234 334574 428854 334658
rect 428234 334338 428266 334574
rect 428502 334338 428586 334574
rect 428822 334338 428854 334574
rect 428234 298894 428854 334338
rect 428234 298658 428266 298894
rect 428502 298658 428586 298894
rect 428822 298658 428854 298894
rect 428234 298574 428854 298658
rect 428234 298338 428266 298574
rect 428502 298338 428586 298574
rect 428822 298338 428854 298574
rect 428234 262894 428854 298338
rect 428234 262658 428266 262894
rect 428502 262658 428586 262894
rect 428822 262658 428854 262894
rect 428234 262574 428854 262658
rect 428234 262338 428266 262574
rect 428502 262338 428586 262574
rect 428822 262338 428854 262574
rect 428234 226894 428854 262338
rect 428234 226658 428266 226894
rect 428502 226658 428586 226894
rect 428822 226658 428854 226894
rect 428234 226574 428854 226658
rect 428234 226338 428266 226574
rect 428502 226338 428586 226574
rect 428822 226338 428854 226574
rect 428234 190894 428854 226338
rect 428234 190658 428266 190894
rect 428502 190658 428586 190894
rect 428822 190658 428854 190894
rect 428234 190574 428854 190658
rect 428234 190338 428266 190574
rect 428502 190338 428586 190574
rect 428822 190338 428854 190574
rect 428234 154894 428854 190338
rect 428234 154658 428266 154894
rect 428502 154658 428586 154894
rect 428822 154658 428854 154894
rect 428234 154574 428854 154658
rect 428234 154338 428266 154574
rect 428502 154338 428586 154574
rect 428822 154338 428854 154574
rect 428234 118894 428854 154338
rect 428234 118658 428266 118894
rect 428502 118658 428586 118894
rect 428822 118658 428854 118894
rect 428234 118574 428854 118658
rect 428234 118338 428266 118574
rect 428502 118338 428586 118574
rect 428822 118338 428854 118574
rect 428234 82894 428854 118338
rect 428234 82658 428266 82894
rect 428502 82658 428586 82894
rect 428822 82658 428854 82894
rect 428234 82574 428854 82658
rect 428234 82338 428266 82574
rect 428502 82338 428586 82574
rect 428822 82338 428854 82574
rect 428234 46894 428854 82338
rect 428234 46658 428266 46894
rect 428502 46658 428586 46894
rect 428822 46658 428854 46894
rect 428234 46574 428854 46658
rect 428234 46338 428266 46574
rect 428502 46338 428586 46574
rect 428822 46338 428854 46574
rect 428234 10894 428854 46338
rect 428234 10658 428266 10894
rect 428502 10658 428586 10894
rect 428822 10658 428854 10894
rect 428234 10574 428854 10658
rect 428234 10338 428266 10574
rect 428502 10338 428586 10574
rect 428822 10338 428854 10574
rect 428234 -4186 428854 10338
rect 430794 705798 431414 705830
rect 430794 705562 430826 705798
rect 431062 705562 431146 705798
rect 431382 705562 431414 705798
rect 430794 705478 431414 705562
rect 430794 705242 430826 705478
rect 431062 705242 431146 705478
rect 431382 705242 431414 705478
rect 430794 669454 431414 705242
rect 430794 669218 430826 669454
rect 431062 669218 431146 669454
rect 431382 669218 431414 669454
rect 430794 669134 431414 669218
rect 430794 668898 430826 669134
rect 431062 668898 431146 669134
rect 431382 668898 431414 669134
rect 430794 633454 431414 668898
rect 430794 633218 430826 633454
rect 431062 633218 431146 633454
rect 431382 633218 431414 633454
rect 430794 633134 431414 633218
rect 430794 632898 430826 633134
rect 431062 632898 431146 633134
rect 431382 632898 431414 633134
rect 430794 597454 431414 632898
rect 430794 597218 430826 597454
rect 431062 597218 431146 597454
rect 431382 597218 431414 597454
rect 430794 597134 431414 597218
rect 430794 596898 430826 597134
rect 431062 596898 431146 597134
rect 431382 596898 431414 597134
rect 430794 561454 431414 596898
rect 430794 561218 430826 561454
rect 431062 561218 431146 561454
rect 431382 561218 431414 561454
rect 430794 561134 431414 561218
rect 430794 560898 430826 561134
rect 431062 560898 431146 561134
rect 431382 560898 431414 561134
rect 430794 525454 431414 560898
rect 430794 525218 430826 525454
rect 431062 525218 431146 525454
rect 431382 525218 431414 525454
rect 430794 525134 431414 525218
rect 430794 524898 430826 525134
rect 431062 524898 431146 525134
rect 431382 524898 431414 525134
rect 430794 489454 431414 524898
rect 430794 489218 430826 489454
rect 431062 489218 431146 489454
rect 431382 489218 431414 489454
rect 430794 489134 431414 489218
rect 430794 488898 430826 489134
rect 431062 488898 431146 489134
rect 431382 488898 431414 489134
rect 430794 453454 431414 488898
rect 430794 453218 430826 453454
rect 431062 453218 431146 453454
rect 431382 453218 431414 453454
rect 430794 453134 431414 453218
rect 430794 452898 430826 453134
rect 431062 452898 431146 453134
rect 431382 452898 431414 453134
rect 430794 417454 431414 452898
rect 430794 417218 430826 417454
rect 431062 417218 431146 417454
rect 431382 417218 431414 417454
rect 430794 417134 431414 417218
rect 430794 416898 430826 417134
rect 431062 416898 431146 417134
rect 431382 416898 431414 417134
rect 430794 381454 431414 416898
rect 430794 381218 430826 381454
rect 431062 381218 431146 381454
rect 431382 381218 431414 381454
rect 430794 381134 431414 381218
rect 430794 380898 430826 381134
rect 431062 380898 431146 381134
rect 431382 380898 431414 381134
rect 430794 345454 431414 380898
rect 430794 345218 430826 345454
rect 431062 345218 431146 345454
rect 431382 345218 431414 345454
rect 430794 345134 431414 345218
rect 430794 344898 430826 345134
rect 431062 344898 431146 345134
rect 431382 344898 431414 345134
rect 430794 309454 431414 344898
rect 430794 309218 430826 309454
rect 431062 309218 431146 309454
rect 431382 309218 431414 309454
rect 430794 309134 431414 309218
rect 430794 308898 430826 309134
rect 431062 308898 431146 309134
rect 431382 308898 431414 309134
rect 430794 273454 431414 308898
rect 430794 273218 430826 273454
rect 431062 273218 431146 273454
rect 431382 273218 431414 273454
rect 430794 273134 431414 273218
rect 430794 272898 430826 273134
rect 431062 272898 431146 273134
rect 431382 272898 431414 273134
rect 430794 237454 431414 272898
rect 430794 237218 430826 237454
rect 431062 237218 431146 237454
rect 431382 237218 431414 237454
rect 430794 237134 431414 237218
rect 430794 236898 430826 237134
rect 431062 236898 431146 237134
rect 431382 236898 431414 237134
rect 430794 201454 431414 236898
rect 430794 201218 430826 201454
rect 431062 201218 431146 201454
rect 431382 201218 431414 201454
rect 430794 201134 431414 201218
rect 430794 200898 430826 201134
rect 431062 200898 431146 201134
rect 431382 200898 431414 201134
rect 430794 165454 431414 200898
rect 430794 165218 430826 165454
rect 431062 165218 431146 165454
rect 431382 165218 431414 165454
rect 430794 165134 431414 165218
rect 430794 164898 430826 165134
rect 431062 164898 431146 165134
rect 431382 164898 431414 165134
rect 430794 129454 431414 164898
rect 430794 129218 430826 129454
rect 431062 129218 431146 129454
rect 431382 129218 431414 129454
rect 430794 129134 431414 129218
rect 430794 128898 430826 129134
rect 431062 128898 431146 129134
rect 431382 128898 431414 129134
rect 430794 93454 431414 128898
rect 430794 93218 430826 93454
rect 431062 93218 431146 93454
rect 431382 93218 431414 93454
rect 430794 93134 431414 93218
rect 430794 92898 430826 93134
rect 431062 92898 431146 93134
rect 431382 92898 431414 93134
rect 430794 57454 431414 92898
rect 430794 57218 430826 57454
rect 431062 57218 431146 57454
rect 431382 57218 431414 57454
rect 430794 57134 431414 57218
rect 430794 56898 430826 57134
rect 431062 56898 431146 57134
rect 431382 56898 431414 57134
rect 430794 21454 431414 56898
rect 430794 21218 430826 21454
rect 431062 21218 431146 21454
rect 431382 21218 431414 21454
rect 430794 21134 431414 21218
rect 430794 20898 430826 21134
rect 431062 20898 431146 21134
rect 431382 20898 431414 21134
rect 430794 -1306 431414 20898
rect 430794 -1542 430826 -1306
rect 431062 -1542 431146 -1306
rect 431382 -1542 431414 -1306
rect 430794 -1626 431414 -1542
rect 430794 -1862 430826 -1626
rect 431062 -1862 431146 -1626
rect 431382 -1862 431414 -1626
rect 430794 -1894 431414 -1862
rect 431954 698614 432574 710042
rect 441954 711558 442574 711590
rect 441954 711322 441986 711558
rect 442222 711322 442306 711558
rect 442542 711322 442574 711558
rect 441954 711238 442574 711322
rect 441954 711002 441986 711238
rect 442222 711002 442306 711238
rect 442542 711002 442574 711238
rect 438234 709638 438854 709670
rect 438234 709402 438266 709638
rect 438502 709402 438586 709638
rect 438822 709402 438854 709638
rect 438234 709318 438854 709402
rect 438234 709082 438266 709318
rect 438502 709082 438586 709318
rect 438822 709082 438854 709318
rect 431954 698378 431986 698614
rect 432222 698378 432306 698614
rect 432542 698378 432574 698614
rect 431954 698294 432574 698378
rect 431954 698058 431986 698294
rect 432222 698058 432306 698294
rect 432542 698058 432574 698294
rect 431954 662614 432574 698058
rect 431954 662378 431986 662614
rect 432222 662378 432306 662614
rect 432542 662378 432574 662614
rect 431954 662294 432574 662378
rect 431954 662058 431986 662294
rect 432222 662058 432306 662294
rect 432542 662058 432574 662294
rect 431954 626614 432574 662058
rect 431954 626378 431986 626614
rect 432222 626378 432306 626614
rect 432542 626378 432574 626614
rect 431954 626294 432574 626378
rect 431954 626058 431986 626294
rect 432222 626058 432306 626294
rect 432542 626058 432574 626294
rect 431954 590614 432574 626058
rect 431954 590378 431986 590614
rect 432222 590378 432306 590614
rect 432542 590378 432574 590614
rect 431954 590294 432574 590378
rect 431954 590058 431986 590294
rect 432222 590058 432306 590294
rect 432542 590058 432574 590294
rect 431954 554614 432574 590058
rect 431954 554378 431986 554614
rect 432222 554378 432306 554614
rect 432542 554378 432574 554614
rect 431954 554294 432574 554378
rect 431954 554058 431986 554294
rect 432222 554058 432306 554294
rect 432542 554058 432574 554294
rect 431954 518614 432574 554058
rect 431954 518378 431986 518614
rect 432222 518378 432306 518614
rect 432542 518378 432574 518614
rect 431954 518294 432574 518378
rect 431954 518058 431986 518294
rect 432222 518058 432306 518294
rect 432542 518058 432574 518294
rect 431954 482614 432574 518058
rect 431954 482378 431986 482614
rect 432222 482378 432306 482614
rect 432542 482378 432574 482614
rect 431954 482294 432574 482378
rect 431954 482058 431986 482294
rect 432222 482058 432306 482294
rect 432542 482058 432574 482294
rect 431954 446614 432574 482058
rect 431954 446378 431986 446614
rect 432222 446378 432306 446614
rect 432542 446378 432574 446614
rect 431954 446294 432574 446378
rect 431954 446058 431986 446294
rect 432222 446058 432306 446294
rect 432542 446058 432574 446294
rect 431954 410614 432574 446058
rect 431954 410378 431986 410614
rect 432222 410378 432306 410614
rect 432542 410378 432574 410614
rect 431954 410294 432574 410378
rect 431954 410058 431986 410294
rect 432222 410058 432306 410294
rect 432542 410058 432574 410294
rect 431954 374614 432574 410058
rect 431954 374378 431986 374614
rect 432222 374378 432306 374614
rect 432542 374378 432574 374614
rect 431954 374294 432574 374378
rect 431954 374058 431986 374294
rect 432222 374058 432306 374294
rect 432542 374058 432574 374294
rect 431954 338614 432574 374058
rect 431954 338378 431986 338614
rect 432222 338378 432306 338614
rect 432542 338378 432574 338614
rect 431954 338294 432574 338378
rect 431954 338058 431986 338294
rect 432222 338058 432306 338294
rect 432542 338058 432574 338294
rect 431954 302614 432574 338058
rect 431954 302378 431986 302614
rect 432222 302378 432306 302614
rect 432542 302378 432574 302614
rect 431954 302294 432574 302378
rect 431954 302058 431986 302294
rect 432222 302058 432306 302294
rect 432542 302058 432574 302294
rect 431954 266614 432574 302058
rect 431954 266378 431986 266614
rect 432222 266378 432306 266614
rect 432542 266378 432574 266614
rect 431954 266294 432574 266378
rect 431954 266058 431986 266294
rect 432222 266058 432306 266294
rect 432542 266058 432574 266294
rect 431954 230614 432574 266058
rect 431954 230378 431986 230614
rect 432222 230378 432306 230614
rect 432542 230378 432574 230614
rect 431954 230294 432574 230378
rect 431954 230058 431986 230294
rect 432222 230058 432306 230294
rect 432542 230058 432574 230294
rect 431954 194614 432574 230058
rect 431954 194378 431986 194614
rect 432222 194378 432306 194614
rect 432542 194378 432574 194614
rect 431954 194294 432574 194378
rect 431954 194058 431986 194294
rect 432222 194058 432306 194294
rect 432542 194058 432574 194294
rect 431954 158614 432574 194058
rect 431954 158378 431986 158614
rect 432222 158378 432306 158614
rect 432542 158378 432574 158614
rect 431954 158294 432574 158378
rect 431954 158058 431986 158294
rect 432222 158058 432306 158294
rect 432542 158058 432574 158294
rect 431954 122614 432574 158058
rect 431954 122378 431986 122614
rect 432222 122378 432306 122614
rect 432542 122378 432574 122614
rect 431954 122294 432574 122378
rect 431954 122058 431986 122294
rect 432222 122058 432306 122294
rect 432542 122058 432574 122294
rect 431954 86614 432574 122058
rect 431954 86378 431986 86614
rect 432222 86378 432306 86614
rect 432542 86378 432574 86614
rect 431954 86294 432574 86378
rect 431954 86058 431986 86294
rect 432222 86058 432306 86294
rect 432542 86058 432574 86294
rect 431954 50614 432574 86058
rect 431954 50378 431986 50614
rect 432222 50378 432306 50614
rect 432542 50378 432574 50614
rect 431954 50294 432574 50378
rect 431954 50058 431986 50294
rect 432222 50058 432306 50294
rect 432542 50058 432574 50294
rect 431954 14614 432574 50058
rect 431954 14378 431986 14614
rect 432222 14378 432306 14614
rect 432542 14378 432574 14614
rect 431954 14294 432574 14378
rect 431954 14058 431986 14294
rect 432222 14058 432306 14294
rect 432542 14058 432574 14294
rect 428234 -4422 428266 -4186
rect 428502 -4422 428586 -4186
rect 428822 -4422 428854 -4186
rect 428234 -4506 428854 -4422
rect 428234 -4742 428266 -4506
rect 428502 -4742 428586 -4506
rect 428822 -4742 428854 -4506
rect 428234 -5734 428854 -4742
rect 421954 -7302 421986 -7066
rect 422222 -7302 422306 -7066
rect 422542 -7302 422574 -7066
rect 421954 -7386 422574 -7302
rect 421954 -7622 421986 -7386
rect 422222 -7622 422306 -7386
rect 422542 -7622 422574 -7386
rect 421954 -7654 422574 -7622
rect 431954 -6106 432574 14058
rect 434514 707718 435134 707750
rect 434514 707482 434546 707718
rect 434782 707482 434866 707718
rect 435102 707482 435134 707718
rect 434514 707398 435134 707482
rect 434514 707162 434546 707398
rect 434782 707162 434866 707398
rect 435102 707162 435134 707398
rect 434514 673174 435134 707162
rect 434514 672938 434546 673174
rect 434782 672938 434866 673174
rect 435102 672938 435134 673174
rect 434514 672854 435134 672938
rect 434514 672618 434546 672854
rect 434782 672618 434866 672854
rect 435102 672618 435134 672854
rect 434514 637174 435134 672618
rect 434514 636938 434546 637174
rect 434782 636938 434866 637174
rect 435102 636938 435134 637174
rect 434514 636854 435134 636938
rect 434514 636618 434546 636854
rect 434782 636618 434866 636854
rect 435102 636618 435134 636854
rect 434514 601174 435134 636618
rect 434514 600938 434546 601174
rect 434782 600938 434866 601174
rect 435102 600938 435134 601174
rect 434514 600854 435134 600938
rect 434514 600618 434546 600854
rect 434782 600618 434866 600854
rect 435102 600618 435134 600854
rect 434514 565174 435134 600618
rect 434514 564938 434546 565174
rect 434782 564938 434866 565174
rect 435102 564938 435134 565174
rect 434514 564854 435134 564938
rect 434514 564618 434546 564854
rect 434782 564618 434866 564854
rect 435102 564618 435134 564854
rect 434514 529174 435134 564618
rect 434514 528938 434546 529174
rect 434782 528938 434866 529174
rect 435102 528938 435134 529174
rect 434514 528854 435134 528938
rect 434514 528618 434546 528854
rect 434782 528618 434866 528854
rect 435102 528618 435134 528854
rect 434514 493174 435134 528618
rect 434514 492938 434546 493174
rect 434782 492938 434866 493174
rect 435102 492938 435134 493174
rect 434514 492854 435134 492938
rect 434514 492618 434546 492854
rect 434782 492618 434866 492854
rect 435102 492618 435134 492854
rect 434514 457174 435134 492618
rect 434514 456938 434546 457174
rect 434782 456938 434866 457174
rect 435102 456938 435134 457174
rect 434514 456854 435134 456938
rect 434514 456618 434546 456854
rect 434782 456618 434866 456854
rect 435102 456618 435134 456854
rect 434514 421174 435134 456618
rect 434514 420938 434546 421174
rect 434782 420938 434866 421174
rect 435102 420938 435134 421174
rect 434514 420854 435134 420938
rect 434514 420618 434546 420854
rect 434782 420618 434866 420854
rect 435102 420618 435134 420854
rect 434514 385174 435134 420618
rect 434514 384938 434546 385174
rect 434782 384938 434866 385174
rect 435102 384938 435134 385174
rect 434514 384854 435134 384938
rect 434514 384618 434546 384854
rect 434782 384618 434866 384854
rect 435102 384618 435134 384854
rect 434514 349174 435134 384618
rect 434514 348938 434546 349174
rect 434782 348938 434866 349174
rect 435102 348938 435134 349174
rect 434514 348854 435134 348938
rect 434514 348618 434546 348854
rect 434782 348618 434866 348854
rect 435102 348618 435134 348854
rect 434514 313174 435134 348618
rect 434514 312938 434546 313174
rect 434782 312938 434866 313174
rect 435102 312938 435134 313174
rect 434514 312854 435134 312938
rect 434514 312618 434546 312854
rect 434782 312618 434866 312854
rect 435102 312618 435134 312854
rect 434514 277174 435134 312618
rect 434514 276938 434546 277174
rect 434782 276938 434866 277174
rect 435102 276938 435134 277174
rect 434514 276854 435134 276938
rect 434514 276618 434546 276854
rect 434782 276618 434866 276854
rect 435102 276618 435134 276854
rect 434514 241174 435134 276618
rect 434514 240938 434546 241174
rect 434782 240938 434866 241174
rect 435102 240938 435134 241174
rect 434514 240854 435134 240938
rect 434514 240618 434546 240854
rect 434782 240618 434866 240854
rect 435102 240618 435134 240854
rect 434514 205174 435134 240618
rect 434514 204938 434546 205174
rect 434782 204938 434866 205174
rect 435102 204938 435134 205174
rect 434514 204854 435134 204938
rect 434514 204618 434546 204854
rect 434782 204618 434866 204854
rect 435102 204618 435134 204854
rect 434514 169174 435134 204618
rect 434514 168938 434546 169174
rect 434782 168938 434866 169174
rect 435102 168938 435134 169174
rect 434514 168854 435134 168938
rect 434514 168618 434546 168854
rect 434782 168618 434866 168854
rect 435102 168618 435134 168854
rect 434514 133174 435134 168618
rect 434514 132938 434546 133174
rect 434782 132938 434866 133174
rect 435102 132938 435134 133174
rect 434514 132854 435134 132938
rect 434514 132618 434546 132854
rect 434782 132618 434866 132854
rect 435102 132618 435134 132854
rect 434514 97174 435134 132618
rect 434514 96938 434546 97174
rect 434782 96938 434866 97174
rect 435102 96938 435134 97174
rect 434514 96854 435134 96938
rect 434514 96618 434546 96854
rect 434782 96618 434866 96854
rect 435102 96618 435134 96854
rect 434514 61174 435134 96618
rect 434514 60938 434546 61174
rect 434782 60938 434866 61174
rect 435102 60938 435134 61174
rect 434514 60854 435134 60938
rect 434514 60618 434546 60854
rect 434782 60618 434866 60854
rect 435102 60618 435134 60854
rect 434514 25174 435134 60618
rect 434514 24938 434546 25174
rect 434782 24938 434866 25174
rect 435102 24938 435134 25174
rect 434514 24854 435134 24938
rect 434514 24618 434546 24854
rect 434782 24618 434866 24854
rect 435102 24618 435134 24854
rect 434514 -3226 435134 24618
rect 434514 -3462 434546 -3226
rect 434782 -3462 434866 -3226
rect 435102 -3462 435134 -3226
rect 434514 -3546 435134 -3462
rect 434514 -3782 434546 -3546
rect 434782 -3782 434866 -3546
rect 435102 -3782 435134 -3546
rect 434514 -3814 435134 -3782
rect 438234 676894 438854 709082
rect 438234 676658 438266 676894
rect 438502 676658 438586 676894
rect 438822 676658 438854 676894
rect 438234 676574 438854 676658
rect 438234 676338 438266 676574
rect 438502 676338 438586 676574
rect 438822 676338 438854 676574
rect 438234 640894 438854 676338
rect 438234 640658 438266 640894
rect 438502 640658 438586 640894
rect 438822 640658 438854 640894
rect 438234 640574 438854 640658
rect 438234 640338 438266 640574
rect 438502 640338 438586 640574
rect 438822 640338 438854 640574
rect 438234 604894 438854 640338
rect 438234 604658 438266 604894
rect 438502 604658 438586 604894
rect 438822 604658 438854 604894
rect 438234 604574 438854 604658
rect 438234 604338 438266 604574
rect 438502 604338 438586 604574
rect 438822 604338 438854 604574
rect 438234 568894 438854 604338
rect 438234 568658 438266 568894
rect 438502 568658 438586 568894
rect 438822 568658 438854 568894
rect 438234 568574 438854 568658
rect 438234 568338 438266 568574
rect 438502 568338 438586 568574
rect 438822 568338 438854 568574
rect 438234 532894 438854 568338
rect 438234 532658 438266 532894
rect 438502 532658 438586 532894
rect 438822 532658 438854 532894
rect 438234 532574 438854 532658
rect 438234 532338 438266 532574
rect 438502 532338 438586 532574
rect 438822 532338 438854 532574
rect 438234 496894 438854 532338
rect 438234 496658 438266 496894
rect 438502 496658 438586 496894
rect 438822 496658 438854 496894
rect 438234 496574 438854 496658
rect 438234 496338 438266 496574
rect 438502 496338 438586 496574
rect 438822 496338 438854 496574
rect 438234 460894 438854 496338
rect 438234 460658 438266 460894
rect 438502 460658 438586 460894
rect 438822 460658 438854 460894
rect 438234 460574 438854 460658
rect 438234 460338 438266 460574
rect 438502 460338 438586 460574
rect 438822 460338 438854 460574
rect 438234 424894 438854 460338
rect 438234 424658 438266 424894
rect 438502 424658 438586 424894
rect 438822 424658 438854 424894
rect 438234 424574 438854 424658
rect 438234 424338 438266 424574
rect 438502 424338 438586 424574
rect 438822 424338 438854 424574
rect 438234 388894 438854 424338
rect 438234 388658 438266 388894
rect 438502 388658 438586 388894
rect 438822 388658 438854 388894
rect 438234 388574 438854 388658
rect 438234 388338 438266 388574
rect 438502 388338 438586 388574
rect 438822 388338 438854 388574
rect 438234 352894 438854 388338
rect 438234 352658 438266 352894
rect 438502 352658 438586 352894
rect 438822 352658 438854 352894
rect 438234 352574 438854 352658
rect 438234 352338 438266 352574
rect 438502 352338 438586 352574
rect 438822 352338 438854 352574
rect 438234 316894 438854 352338
rect 438234 316658 438266 316894
rect 438502 316658 438586 316894
rect 438822 316658 438854 316894
rect 438234 316574 438854 316658
rect 438234 316338 438266 316574
rect 438502 316338 438586 316574
rect 438822 316338 438854 316574
rect 438234 280894 438854 316338
rect 438234 280658 438266 280894
rect 438502 280658 438586 280894
rect 438822 280658 438854 280894
rect 438234 280574 438854 280658
rect 438234 280338 438266 280574
rect 438502 280338 438586 280574
rect 438822 280338 438854 280574
rect 438234 244894 438854 280338
rect 438234 244658 438266 244894
rect 438502 244658 438586 244894
rect 438822 244658 438854 244894
rect 438234 244574 438854 244658
rect 438234 244338 438266 244574
rect 438502 244338 438586 244574
rect 438822 244338 438854 244574
rect 438234 208894 438854 244338
rect 438234 208658 438266 208894
rect 438502 208658 438586 208894
rect 438822 208658 438854 208894
rect 438234 208574 438854 208658
rect 438234 208338 438266 208574
rect 438502 208338 438586 208574
rect 438822 208338 438854 208574
rect 438234 172894 438854 208338
rect 438234 172658 438266 172894
rect 438502 172658 438586 172894
rect 438822 172658 438854 172894
rect 438234 172574 438854 172658
rect 438234 172338 438266 172574
rect 438502 172338 438586 172574
rect 438822 172338 438854 172574
rect 438234 136894 438854 172338
rect 438234 136658 438266 136894
rect 438502 136658 438586 136894
rect 438822 136658 438854 136894
rect 438234 136574 438854 136658
rect 438234 136338 438266 136574
rect 438502 136338 438586 136574
rect 438822 136338 438854 136574
rect 438234 100894 438854 136338
rect 438234 100658 438266 100894
rect 438502 100658 438586 100894
rect 438822 100658 438854 100894
rect 438234 100574 438854 100658
rect 438234 100338 438266 100574
rect 438502 100338 438586 100574
rect 438822 100338 438854 100574
rect 438234 64894 438854 100338
rect 438234 64658 438266 64894
rect 438502 64658 438586 64894
rect 438822 64658 438854 64894
rect 438234 64574 438854 64658
rect 438234 64338 438266 64574
rect 438502 64338 438586 64574
rect 438822 64338 438854 64574
rect 438234 28894 438854 64338
rect 438234 28658 438266 28894
rect 438502 28658 438586 28894
rect 438822 28658 438854 28894
rect 438234 28574 438854 28658
rect 438234 28338 438266 28574
rect 438502 28338 438586 28574
rect 438822 28338 438854 28574
rect 438234 -5146 438854 28338
rect 440794 704838 441414 705830
rect 440794 704602 440826 704838
rect 441062 704602 441146 704838
rect 441382 704602 441414 704838
rect 440794 704518 441414 704602
rect 440794 704282 440826 704518
rect 441062 704282 441146 704518
rect 441382 704282 441414 704518
rect 440794 687454 441414 704282
rect 440794 687218 440826 687454
rect 441062 687218 441146 687454
rect 441382 687218 441414 687454
rect 440794 687134 441414 687218
rect 440794 686898 440826 687134
rect 441062 686898 441146 687134
rect 441382 686898 441414 687134
rect 440794 651454 441414 686898
rect 440794 651218 440826 651454
rect 441062 651218 441146 651454
rect 441382 651218 441414 651454
rect 440794 651134 441414 651218
rect 440794 650898 440826 651134
rect 441062 650898 441146 651134
rect 441382 650898 441414 651134
rect 440794 615454 441414 650898
rect 440794 615218 440826 615454
rect 441062 615218 441146 615454
rect 441382 615218 441414 615454
rect 440794 615134 441414 615218
rect 440794 614898 440826 615134
rect 441062 614898 441146 615134
rect 441382 614898 441414 615134
rect 440794 579454 441414 614898
rect 440794 579218 440826 579454
rect 441062 579218 441146 579454
rect 441382 579218 441414 579454
rect 440794 579134 441414 579218
rect 440794 578898 440826 579134
rect 441062 578898 441146 579134
rect 441382 578898 441414 579134
rect 440794 543454 441414 578898
rect 440794 543218 440826 543454
rect 441062 543218 441146 543454
rect 441382 543218 441414 543454
rect 440794 543134 441414 543218
rect 440794 542898 440826 543134
rect 441062 542898 441146 543134
rect 441382 542898 441414 543134
rect 440794 507454 441414 542898
rect 440794 507218 440826 507454
rect 441062 507218 441146 507454
rect 441382 507218 441414 507454
rect 440794 507134 441414 507218
rect 440794 506898 440826 507134
rect 441062 506898 441146 507134
rect 441382 506898 441414 507134
rect 440794 471454 441414 506898
rect 440794 471218 440826 471454
rect 441062 471218 441146 471454
rect 441382 471218 441414 471454
rect 440794 471134 441414 471218
rect 440794 470898 440826 471134
rect 441062 470898 441146 471134
rect 441382 470898 441414 471134
rect 440794 435454 441414 470898
rect 440794 435218 440826 435454
rect 441062 435218 441146 435454
rect 441382 435218 441414 435454
rect 440794 435134 441414 435218
rect 440794 434898 440826 435134
rect 441062 434898 441146 435134
rect 441382 434898 441414 435134
rect 440794 399454 441414 434898
rect 440794 399218 440826 399454
rect 441062 399218 441146 399454
rect 441382 399218 441414 399454
rect 440794 399134 441414 399218
rect 440794 398898 440826 399134
rect 441062 398898 441146 399134
rect 441382 398898 441414 399134
rect 440794 363454 441414 398898
rect 440794 363218 440826 363454
rect 441062 363218 441146 363454
rect 441382 363218 441414 363454
rect 440794 363134 441414 363218
rect 440794 362898 440826 363134
rect 441062 362898 441146 363134
rect 441382 362898 441414 363134
rect 440794 327454 441414 362898
rect 440794 327218 440826 327454
rect 441062 327218 441146 327454
rect 441382 327218 441414 327454
rect 440794 327134 441414 327218
rect 440794 326898 440826 327134
rect 441062 326898 441146 327134
rect 441382 326898 441414 327134
rect 440794 291454 441414 326898
rect 440794 291218 440826 291454
rect 441062 291218 441146 291454
rect 441382 291218 441414 291454
rect 440794 291134 441414 291218
rect 440794 290898 440826 291134
rect 441062 290898 441146 291134
rect 441382 290898 441414 291134
rect 440794 255454 441414 290898
rect 440794 255218 440826 255454
rect 441062 255218 441146 255454
rect 441382 255218 441414 255454
rect 440794 255134 441414 255218
rect 440794 254898 440826 255134
rect 441062 254898 441146 255134
rect 441382 254898 441414 255134
rect 440794 219454 441414 254898
rect 440794 219218 440826 219454
rect 441062 219218 441146 219454
rect 441382 219218 441414 219454
rect 440794 219134 441414 219218
rect 440794 218898 440826 219134
rect 441062 218898 441146 219134
rect 441382 218898 441414 219134
rect 440794 183454 441414 218898
rect 440794 183218 440826 183454
rect 441062 183218 441146 183454
rect 441382 183218 441414 183454
rect 440794 183134 441414 183218
rect 440794 182898 440826 183134
rect 441062 182898 441146 183134
rect 441382 182898 441414 183134
rect 440794 147454 441414 182898
rect 440794 147218 440826 147454
rect 441062 147218 441146 147454
rect 441382 147218 441414 147454
rect 440794 147134 441414 147218
rect 440794 146898 440826 147134
rect 441062 146898 441146 147134
rect 441382 146898 441414 147134
rect 440794 111454 441414 146898
rect 440794 111218 440826 111454
rect 441062 111218 441146 111454
rect 441382 111218 441414 111454
rect 440794 111134 441414 111218
rect 440794 110898 440826 111134
rect 441062 110898 441146 111134
rect 441382 110898 441414 111134
rect 440794 75454 441414 110898
rect 440794 75218 440826 75454
rect 441062 75218 441146 75454
rect 441382 75218 441414 75454
rect 440794 75134 441414 75218
rect 440794 74898 440826 75134
rect 441062 74898 441146 75134
rect 441382 74898 441414 75134
rect 440794 39454 441414 74898
rect 440794 39218 440826 39454
rect 441062 39218 441146 39454
rect 441382 39218 441414 39454
rect 440794 39134 441414 39218
rect 440794 38898 440826 39134
rect 441062 38898 441146 39134
rect 441382 38898 441414 39134
rect 440794 3454 441414 38898
rect 440794 3218 440826 3454
rect 441062 3218 441146 3454
rect 441382 3218 441414 3454
rect 440794 3134 441414 3218
rect 440794 2898 440826 3134
rect 441062 2898 441146 3134
rect 441382 2898 441414 3134
rect 440794 -346 441414 2898
rect 440794 -582 440826 -346
rect 441062 -582 441146 -346
rect 441382 -582 441414 -346
rect 440794 -666 441414 -582
rect 440794 -902 440826 -666
rect 441062 -902 441146 -666
rect 441382 -902 441414 -666
rect 440794 -1894 441414 -902
rect 441954 680614 442574 711002
rect 451954 710598 452574 711590
rect 451954 710362 451986 710598
rect 452222 710362 452306 710598
rect 452542 710362 452574 710598
rect 451954 710278 452574 710362
rect 451954 710042 451986 710278
rect 452222 710042 452306 710278
rect 452542 710042 452574 710278
rect 448234 708678 448854 709670
rect 448234 708442 448266 708678
rect 448502 708442 448586 708678
rect 448822 708442 448854 708678
rect 448234 708358 448854 708442
rect 448234 708122 448266 708358
rect 448502 708122 448586 708358
rect 448822 708122 448854 708358
rect 441954 680378 441986 680614
rect 442222 680378 442306 680614
rect 442542 680378 442574 680614
rect 441954 680294 442574 680378
rect 441954 680058 441986 680294
rect 442222 680058 442306 680294
rect 442542 680058 442574 680294
rect 441954 644614 442574 680058
rect 441954 644378 441986 644614
rect 442222 644378 442306 644614
rect 442542 644378 442574 644614
rect 441954 644294 442574 644378
rect 441954 644058 441986 644294
rect 442222 644058 442306 644294
rect 442542 644058 442574 644294
rect 441954 608614 442574 644058
rect 441954 608378 441986 608614
rect 442222 608378 442306 608614
rect 442542 608378 442574 608614
rect 441954 608294 442574 608378
rect 441954 608058 441986 608294
rect 442222 608058 442306 608294
rect 442542 608058 442574 608294
rect 441954 572614 442574 608058
rect 441954 572378 441986 572614
rect 442222 572378 442306 572614
rect 442542 572378 442574 572614
rect 441954 572294 442574 572378
rect 441954 572058 441986 572294
rect 442222 572058 442306 572294
rect 442542 572058 442574 572294
rect 441954 536614 442574 572058
rect 441954 536378 441986 536614
rect 442222 536378 442306 536614
rect 442542 536378 442574 536614
rect 441954 536294 442574 536378
rect 441954 536058 441986 536294
rect 442222 536058 442306 536294
rect 442542 536058 442574 536294
rect 441954 500614 442574 536058
rect 441954 500378 441986 500614
rect 442222 500378 442306 500614
rect 442542 500378 442574 500614
rect 441954 500294 442574 500378
rect 441954 500058 441986 500294
rect 442222 500058 442306 500294
rect 442542 500058 442574 500294
rect 441954 464614 442574 500058
rect 441954 464378 441986 464614
rect 442222 464378 442306 464614
rect 442542 464378 442574 464614
rect 441954 464294 442574 464378
rect 441954 464058 441986 464294
rect 442222 464058 442306 464294
rect 442542 464058 442574 464294
rect 441954 428614 442574 464058
rect 441954 428378 441986 428614
rect 442222 428378 442306 428614
rect 442542 428378 442574 428614
rect 441954 428294 442574 428378
rect 441954 428058 441986 428294
rect 442222 428058 442306 428294
rect 442542 428058 442574 428294
rect 441954 392614 442574 428058
rect 441954 392378 441986 392614
rect 442222 392378 442306 392614
rect 442542 392378 442574 392614
rect 441954 392294 442574 392378
rect 441954 392058 441986 392294
rect 442222 392058 442306 392294
rect 442542 392058 442574 392294
rect 441954 356614 442574 392058
rect 441954 356378 441986 356614
rect 442222 356378 442306 356614
rect 442542 356378 442574 356614
rect 441954 356294 442574 356378
rect 441954 356058 441986 356294
rect 442222 356058 442306 356294
rect 442542 356058 442574 356294
rect 441954 320614 442574 356058
rect 441954 320378 441986 320614
rect 442222 320378 442306 320614
rect 442542 320378 442574 320614
rect 441954 320294 442574 320378
rect 441954 320058 441986 320294
rect 442222 320058 442306 320294
rect 442542 320058 442574 320294
rect 441954 284614 442574 320058
rect 441954 284378 441986 284614
rect 442222 284378 442306 284614
rect 442542 284378 442574 284614
rect 441954 284294 442574 284378
rect 441954 284058 441986 284294
rect 442222 284058 442306 284294
rect 442542 284058 442574 284294
rect 441954 248614 442574 284058
rect 441954 248378 441986 248614
rect 442222 248378 442306 248614
rect 442542 248378 442574 248614
rect 441954 248294 442574 248378
rect 441954 248058 441986 248294
rect 442222 248058 442306 248294
rect 442542 248058 442574 248294
rect 441954 212614 442574 248058
rect 441954 212378 441986 212614
rect 442222 212378 442306 212614
rect 442542 212378 442574 212614
rect 441954 212294 442574 212378
rect 441954 212058 441986 212294
rect 442222 212058 442306 212294
rect 442542 212058 442574 212294
rect 441954 176614 442574 212058
rect 441954 176378 441986 176614
rect 442222 176378 442306 176614
rect 442542 176378 442574 176614
rect 441954 176294 442574 176378
rect 441954 176058 441986 176294
rect 442222 176058 442306 176294
rect 442542 176058 442574 176294
rect 441954 140614 442574 176058
rect 441954 140378 441986 140614
rect 442222 140378 442306 140614
rect 442542 140378 442574 140614
rect 441954 140294 442574 140378
rect 441954 140058 441986 140294
rect 442222 140058 442306 140294
rect 442542 140058 442574 140294
rect 441954 104614 442574 140058
rect 441954 104378 441986 104614
rect 442222 104378 442306 104614
rect 442542 104378 442574 104614
rect 441954 104294 442574 104378
rect 441954 104058 441986 104294
rect 442222 104058 442306 104294
rect 442542 104058 442574 104294
rect 441954 68614 442574 104058
rect 441954 68378 441986 68614
rect 442222 68378 442306 68614
rect 442542 68378 442574 68614
rect 441954 68294 442574 68378
rect 441954 68058 441986 68294
rect 442222 68058 442306 68294
rect 442542 68058 442574 68294
rect 441954 32614 442574 68058
rect 441954 32378 441986 32614
rect 442222 32378 442306 32614
rect 442542 32378 442574 32614
rect 441954 32294 442574 32378
rect 441954 32058 441986 32294
rect 442222 32058 442306 32294
rect 442542 32058 442574 32294
rect 438234 -5382 438266 -5146
rect 438502 -5382 438586 -5146
rect 438822 -5382 438854 -5146
rect 438234 -5466 438854 -5382
rect 438234 -5702 438266 -5466
rect 438502 -5702 438586 -5466
rect 438822 -5702 438854 -5466
rect 438234 -5734 438854 -5702
rect 431954 -6342 431986 -6106
rect 432222 -6342 432306 -6106
rect 432542 -6342 432574 -6106
rect 431954 -6426 432574 -6342
rect 431954 -6662 431986 -6426
rect 432222 -6662 432306 -6426
rect 432542 -6662 432574 -6426
rect 431954 -7654 432574 -6662
rect 441954 -7066 442574 32058
rect 444514 706758 445134 707750
rect 444514 706522 444546 706758
rect 444782 706522 444866 706758
rect 445102 706522 445134 706758
rect 444514 706438 445134 706522
rect 444514 706202 444546 706438
rect 444782 706202 444866 706438
rect 445102 706202 445134 706438
rect 444514 691174 445134 706202
rect 444514 690938 444546 691174
rect 444782 690938 444866 691174
rect 445102 690938 445134 691174
rect 444514 690854 445134 690938
rect 444514 690618 444546 690854
rect 444782 690618 444866 690854
rect 445102 690618 445134 690854
rect 444514 655174 445134 690618
rect 444514 654938 444546 655174
rect 444782 654938 444866 655174
rect 445102 654938 445134 655174
rect 444514 654854 445134 654938
rect 444514 654618 444546 654854
rect 444782 654618 444866 654854
rect 445102 654618 445134 654854
rect 444514 619174 445134 654618
rect 444514 618938 444546 619174
rect 444782 618938 444866 619174
rect 445102 618938 445134 619174
rect 444514 618854 445134 618938
rect 444514 618618 444546 618854
rect 444782 618618 444866 618854
rect 445102 618618 445134 618854
rect 444514 583174 445134 618618
rect 444514 582938 444546 583174
rect 444782 582938 444866 583174
rect 445102 582938 445134 583174
rect 444514 582854 445134 582938
rect 444514 582618 444546 582854
rect 444782 582618 444866 582854
rect 445102 582618 445134 582854
rect 444514 547174 445134 582618
rect 444514 546938 444546 547174
rect 444782 546938 444866 547174
rect 445102 546938 445134 547174
rect 444514 546854 445134 546938
rect 444514 546618 444546 546854
rect 444782 546618 444866 546854
rect 445102 546618 445134 546854
rect 444514 511174 445134 546618
rect 444514 510938 444546 511174
rect 444782 510938 444866 511174
rect 445102 510938 445134 511174
rect 444514 510854 445134 510938
rect 444514 510618 444546 510854
rect 444782 510618 444866 510854
rect 445102 510618 445134 510854
rect 444514 475174 445134 510618
rect 444514 474938 444546 475174
rect 444782 474938 444866 475174
rect 445102 474938 445134 475174
rect 444514 474854 445134 474938
rect 444514 474618 444546 474854
rect 444782 474618 444866 474854
rect 445102 474618 445134 474854
rect 444514 439174 445134 474618
rect 444514 438938 444546 439174
rect 444782 438938 444866 439174
rect 445102 438938 445134 439174
rect 444514 438854 445134 438938
rect 444514 438618 444546 438854
rect 444782 438618 444866 438854
rect 445102 438618 445134 438854
rect 444514 403174 445134 438618
rect 444514 402938 444546 403174
rect 444782 402938 444866 403174
rect 445102 402938 445134 403174
rect 444514 402854 445134 402938
rect 444514 402618 444546 402854
rect 444782 402618 444866 402854
rect 445102 402618 445134 402854
rect 444514 367174 445134 402618
rect 444514 366938 444546 367174
rect 444782 366938 444866 367174
rect 445102 366938 445134 367174
rect 444514 366854 445134 366938
rect 444514 366618 444546 366854
rect 444782 366618 444866 366854
rect 445102 366618 445134 366854
rect 444514 331174 445134 366618
rect 444514 330938 444546 331174
rect 444782 330938 444866 331174
rect 445102 330938 445134 331174
rect 444514 330854 445134 330938
rect 444514 330618 444546 330854
rect 444782 330618 444866 330854
rect 445102 330618 445134 330854
rect 444514 295174 445134 330618
rect 444514 294938 444546 295174
rect 444782 294938 444866 295174
rect 445102 294938 445134 295174
rect 444514 294854 445134 294938
rect 444514 294618 444546 294854
rect 444782 294618 444866 294854
rect 445102 294618 445134 294854
rect 444514 259174 445134 294618
rect 444514 258938 444546 259174
rect 444782 258938 444866 259174
rect 445102 258938 445134 259174
rect 444514 258854 445134 258938
rect 444514 258618 444546 258854
rect 444782 258618 444866 258854
rect 445102 258618 445134 258854
rect 444514 223174 445134 258618
rect 444514 222938 444546 223174
rect 444782 222938 444866 223174
rect 445102 222938 445134 223174
rect 444514 222854 445134 222938
rect 444514 222618 444546 222854
rect 444782 222618 444866 222854
rect 445102 222618 445134 222854
rect 444514 187174 445134 222618
rect 444514 186938 444546 187174
rect 444782 186938 444866 187174
rect 445102 186938 445134 187174
rect 444514 186854 445134 186938
rect 444514 186618 444546 186854
rect 444782 186618 444866 186854
rect 445102 186618 445134 186854
rect 444514 151174 445134 186618
rect 444514 150938 444546 151174
rect 444782 150938 444866 151174
rect 445102 150938 445134 151174
rect 444514 150854 445134 150938
rect 444514 150618 444546 150854
rect 444782 150618 444866 150854
rect 445102 150618 445134 150854
rect 444514 115174 445134 150618
rect 444514 114938 444546 115174
rect 444782 114938 444866 115174
rect 445102 114938 445134 115174
rect 444514 114854 445134 114938
rect 444514 114618 444546 114854
rect 444782 114618 444866 114854
rect 445102 114618 445134 114854
rect 444514 79174 445134 114618
rect 444514 78938 444546 79174
rect 444782 78938 444866 79174
rect 445102 78938 445134 79174
rect 444514 78854 445134 78938
rect 444514 78618 444546 78854
rect 444782 78618 444866 78854
rect 445102 78618 445134 78854
rect 444514 43174 445134 78618
rect 444514 42938 444546 43174
rect 444782 42938 444866 43174
rect 445102 42938 445134 43174
rect 444514 42854 445134 42938
rect 444514 42618 444546 42854
rect 444782 42618 444866 42854
rect 445102 42618 445134 42854
rect 444514 7174 445134 42618
rect 444514 6938 444546 7174
rect 444782 6938 444866 7174
rect 445102 6938 445134 7174
rect 444514 6854 445134 6938
rect 444514 6618 444546 6854
rect 444782 6618 444866 6854
rect 445102 6618 445134 6854
rect 444514 -2266 445134 6618
rect 444514 -2502 444546 -2266
rect 444782 -2502 444866 -2266
rect 445102 -2502 445134 -2266
rect 444514 -2586 445134 -2502
rect 444514 -2822 444546 -2586
rect 444782 -2822 444866 -2586
rect 445102 -2822 445134 -2586
rect 444514 -3814 445134 -2822
rect 448234 694894 448854 708122
rect 448234 694658 448266 694894
rect 448502 694658 448586 694894
rect 448822 694658 448854 694894
rect 448234 694574 448854 694658
rect 448234 694338 448266 694574
rect 448502 694338 448586 694574
rect 448822 694338 448854 694574
rect 448234 658894 448854 694338
rect 448234 658658 448266 658894
rect 448502 658658 448586 658894
rect 448822 658658 448854 658894
rect 448234 658574 448854 658658
rect 448234 658338 448266 658574
rect 448502 658338 448586 658574
rect 448822 658338 448854 658574
rect 448234 622894 448854 658338
rect 448234 622658 448266 622894
rect 448502 622658 448586 622894
rect 448822 622658 448854 622894
rect 448234 622574 448854 622658
rect 448234 622338 448266 622574
rect 448502 622338 448586 622574
rect 448822 622338 448854 622574
rect 448234 586894 448854 622338
rect 448234 586658 448266 586894
rect 448502 586658 448586 586894
rect 448822 586658 448854 586894
rect 448234 586574 448854 586658
rect 448234 586338 448266 586574
rect 448502 586338 448586 586574
rect 448822 586338 448854 586574
rect 448234 550894 448854 586338
rect 448234 550658 448266 550894
rect 448502 550658 448586 550894
rect 448822 550658 448854 550894
rect 448234 550574 448854 550658
rect 448234 550338 448266 550574
rect 448502 550338 448586 550574
rect 448822 550338 448854 550574
rect 448234 514894 448854 550338
rect 448234 514658 448266 514894
rect 448502 514658 448586 514894
rect 448822 514658 448854 514894
rect 448234 514574 448854 514658
rect 448234 514338 448266 514574
rect 448502 514338 448586 514574
rect 448822 514338 448854 514574
rect 448234 478894 448854 514338
rect 448234 478658 448266 478894
rect 448502 478658 448586 478894
rect 448822 478658 448854 478894
rect 448234 478574 448854 478658
rect 448234 478338 448266 478574
rect 448502 478338 448586 478574
rect 448822 478338 448854 478574
rect 448234 442894 448854 478338
rect 448234 442658 448266 442894
rect 448502 442658 448586 442894
rect 448822 442658 448854 442894
rect 448234 442574 448854 442658
rect 448234 442338 448266 442574
rect 448502 442338 448586 442574
rect 448822 442338 448854 442574
rect 448234 406894 448854 442338
rect 448234 406658 448266 406894
rect 448502 406658 448586 406894
rect 448822 406658 448854 406894
rect 448234 406574 448854 406658
rect 448234 406338 448266 406574
rect 448502 406338 448586 406574
rect 448822 406338 448854 406574
rect 448234 370894 448854 406338
rect 448234 370658 448266 370894
rect 448502 370658 448586 370894
rect 448822 370658 448854 370894
rect 448234 370574 448854 370658
rect 448234 370338 448266 370574
rect 448502 370338 448586 370574
rect 448822 370338 448854 370574
rect 448234 334894 448854 370338
rect 448234 334658 448266 334894
rect 448502 334658 448586 334894
rect 448822 334658 448854 334894
rect 448234 334574 448854 334658
rect 448234 334338 448266 334574
rect 448502 334338 448586 334574
rect 448822 334338 448854 334574
rect 448234 298894 448854 334338
rect 448234 298658 448266 298894
rect 448502 298658 448586 298894
rect 448822 298658 448854 298894
rect 448234 298574 448854 298658
rect 448234 298338 448266 298574
rect 448502 298338 448586 298574
rect 448822 298338 448854 298574
rect 448234 262894 448854 298338
rect 448234 262658 448266 262894
rect 448502 262658 448586 262894
rect 448822 262658 448854 262894
rect 448234 262574 448854 262658
rect 448234 262338 448266 262574
rect 448502 262338 448586 262574
rect 448822 262338 448854 262574
rect 448234 226894 448854 262338
rect 448234 226658 448266 226894
rect 448502 226658 448586 226894
rect 448822 226658 448854 226894
rect 448234 226574 448854 226658
rect 448234 226338 448266 226574
rect 448502 226338 448586 226574
rect 448822 226338 448854 226574
rect 448234 190894 448854 226338
rect 448234 190658 448266 190894
rect 448502 190658 448586 190894
rect 448822 190658 448854 190894
rect 448234 190574 448854 190658
rect 448234 190338 448266 190574
rect 448502 190338 448586 190574
rect 448822 190338 448854 190574
rect 448234 154894 448854 190338
rect 448234 154658 448266 154894
rect 448502 154658 448586 154894
rect 448822 154658 448854 154894
rect 448234 154574 448854 154658
rect 448234 154338 448266 154574
rect 448502 154338 448586 154574
rect 448822 154338 448854 154574
rect 448234 118894 448854 154338
rect 448234 118658 448266 118894
rect 448502 118658 448586 118894
rect 448822 118658 448854 118894
rect 448234 118574 448854 118658
rect 448234 118338 448266 118574
rect 448502 118338 448586 118574
rect 448822 118338 448854 118574
rect 448234 82894 448854 118338
rect 448234 82658 448266 82894
rect 448502 82658 448586 82894
rect 448822 82658 448854 82894
rect 448234 82574 448854 82658
rect 448234 82338 448266 82574
rect 448502 82338 448586 82574
rect 448822 82338 448854 82574
rect 448234 46894 448854 82338
rect 448234 46658 448266 46894
rect 448502 46658 448586 46894
rect 448822 46658 448854 46894
rect 448234 46574 448854 46658
rect 448234 46338 448266 46574
rect 448502 46338 448586 46574
rect 448822 46338 448854 46574
rect 448234 10894 448854 46338
rect 448234 10658 448266 10894
rect 448502 10658 448586 10894
rect 448822 10658 448854 10894
rect 448234 10574 448854 10658
rect 448234 10338 448266 10574
rect 448502 10338 448586 10574
rect 448822 10338 448854 10574
rect 448234 -4186 448854 10338
rect 450794 705798 451414 705830
rect 450794 705562 450826 705798
rect 451062 705562 451146 705798
rect 451382 705562 451414 705798
rect 450794 705478 451414 705562
rect 450794 705242 450826 705478
rect 451062 705242 451146 705478
rect 451382 705242 451414 705478
rect 450794 669454 451414 705242
rect 450794 669218 450826 669454
rect 451062 669218 451146 669454
rect 451382 669218 451414 669454
rect 450794 669134 451414 669218
rect 450794 668898 450826 669134
rect 451062 668898 451146 669134
rect 451382 668898 451414 669134
rect 450794 633454 451414 668898
rect 450794 633218 450826 633454
rect 451062 633218 451146 633454
rect 451382 633218 451414 633454
rect 450794 633134 451414 633218
rect 450794 632898 450826 633134
rect 451062 632898 451146 633134
rect 451382 632898 451414 633134
rect 450794 597454 451414 632898
rect 450794 597218 450826 597454
rect 451062 597218 451146 597454
rect 451382 597218 451414 597454
rect 450794 597134 451414 597218
rect 450794 596898 450826 597134
rect 451062 596898 451146 597134
rect 451382 596898 451414 597134
rect 450794 561454 451414 596898
rect 450794 561218 450826 561454
rect 451062 561218 451146 561454
rect 451382 561218 451414 561454
rect 450794 561134 451414 561218
rect 450794 560898 450826 561134
rect 451062 560898 451146 561134
rect 451382 560898 451414 561134
rect 450794 525454 451414 560898
rect 450794 525218 450826 525454
rect 451062 525218 451146 525454
rect 451382 525218 451414 525454
rect 450794 525134 451414 525218
rect 450794 524898 450826 525134
rect 451062 524898 451146 525134
rect 451382 524898 451414 525134
rect 450794 489454 451414 524898
rect 450794 489218 450826 489454
rect 451062 489218 451146 489454
rect 451382 489218 451414 489454
rect 450794 489134 451414 489218
rect 450794 488898 450826 489134
rect 451062 488898 451146 489134
rect 451382 488898 451414 489134
rect 450794 453454 451414 488898
rect 450794 453218 450826 453454
rect 451062 453218 451146 453454
rect 451382 453218 451414 453454
rect 450794 453134 451414 453218
rect 450794 452898 450826 453134
rect 451062 452898 451146 453134
rect 451382 452898 451414 453134
rect 450794 417454 451414 452898
rect 450794 417218 450826 417454
rect 451062 417218 451146 417454
rect 451382 417218 451414 417454
rect 450794 417134 451414 417218
rect 450794 416898 450826 417134
rect 451062 416898 451146 417134
rect 451382 416898 451414 417134
rect 450794 381454 451414 416898
rect 450794 381218 450826 381454
rect 451062 381218 451146 381454
rect 451382 381218 451414 381454
rect 450794 381134 451414 381218
rect 450794 380898 450826 381134
rect 451062 380898 451146 381134
rect 451382 380898 451414 381134
rect 450794 345454 451414 380898
rect 450794 345218 450826 345454
rect 451062 345218 451146 345454
rect 451382 345218 451414 345454
rect 450794 345134 451414 345218
rect 450794 344898 450826 345134
rect 451062 344898 451146 345134
rect 451382 344898 451414 345134
rect 450794 309454 451414 344898
rect 450794 309218 450826 309454
rect 451062 309218 451146 309454
rect 451382 309218 451414 309454
rect 450794 309134 451414 309218
rect 450794 308898 450826 309134
rect 451062 308898 451146 309134
rect 451382 308898 451414 309134
rect 450794 273454 451414 308898
rect 450794 273218 450826 273454
rect 451062 273218 451146 273454
rect 451382 273218 451414 273454
rect 450794 273134 451414 273218
rect 450794 272898 450826 273134
rect 451062 272898 451146 273134
rect 451382 272898 451414 273134
rect 450794 237454 451414 272898
rect 450794 237218 450826 237454
rect 451062 237218 451146 237454
rect 451382 237218 451414 237454
rect 450794 237134 451414 237218
rect 450794 236898 450826 237134
rect 451062 236898 451146 237134
rect 451382 236898 451414 237134
rect 450794 201454 451414 236898
rect 450794 201218 450826 201454
rect 451062 201218 451146 201454
rect 451382 201218 451414 201454
rect 450794 201134 451414 201218
rect 450794 200898 450826 201134
rect 451062 200898 451146 201134
rect 451382 200898 451414 201134
rect 450794 165454 451414 200898
rect 450794 165218 450826 165454
rect 451062 165218 451146 165454
rect 451382 165218 451414 165454
rect 450794 165134 451414 165218
rect 450794 164898 450826 165134
rect 451062 164898 451146 165134
rect 451382 164898 451414 165134
rect 450794 129454 451414 164898
rect 450794 129218 450826 129454
rect 451062 129218 451146 129454
rect 451382 129218 451414 129454
rect 450794 129134 451414 129218
rect 450794 128898 450826 129134
rect 451062 128898 451146 129134
rect 451382 128898 451414 129134
rect 450794 93454 451414 128898
rect 450794 93218 450826 93454
rect 451062 93218 451146 93454
rect 451382 93218 451414 93454
rect 450794 93134 451414 93218
rect 450794 92898 450826 93134
rect 451062 92898 451146 93134
rect 451382 92898 451414 93134
rect 450794 57454 451414 92898
rect 450794 57218 450826 57454
rect 451062 57218 451146 57454
rect 451382 57218 451414 57454
rect 450794 57134 451414 57218
rect 450794 56898 450826 57134
rect 451062 56898 451146 57134
rect 451382 56898 451414 57134
rect 450794 21454 451414 56898
rect 450794 21218 450826 21454
rect 451062 21218 451146 21454
rect 451382 21218 451414 21454
rect 450794 21134 451414 21218
rect 450794 20898 450826 21134
rect 451062 20898 451146 21134
rect 451382 20898 451414 21134
rect 450794 -1306 451414 20898
rect 450794 -1542 450826 -1306
rect 451062 -1542 451146 -1306
rect 451382 -1542 451414 -1306
rect 450794 -1626 451414 -1542
rect 450794 -1862 450826 -1626
rect 451062 -1862 451146 -1626
rect 451382 -1862 451414 -1626
rect 450794 -1894 451414 -1862
rect 451954 698614 452574 710042
rect 461954 711558 462574 711590
rect 461954 711322 461986 711558
rect 462222 711322 462306 711558
rect 462542 711322 462574 711558
rect 461954 711238 462574 711322
rect 461954 711002 461986 711238
rect 462222 711002 462306 711238
rect 462542 711002 462574 711238
rect 458234 709638 458854 709670
rect 458234 709402 458266 709638
rect 458502 709402 458586 709638
rect 458822 709402 458854 709638
rect 458234 709318 458854 709402
rect 458234 709082 458266 709318
rect 458502 709082 458586 709318
rect 458822 709082 458854 709318
rect 451954 698378 451986 698614
rect 452222 698378 452306 698614
rect 452542 698378 452574 698614
rect 451954 698294 452574 698378
rect 451954 698058 451986 698294
rect 452222 698058 452306 698294
rect 452542 698058 452574 698294
rect 451954 662614 452574 698058
rect 451954 662378 451986 662614
rect 452222 662378 452306 662614
rect 452542 662378 452574 662614
rect 451954 662294 452574 662378
rect 451954 662058 451986 662294
rect 452222 662058 452306 662294
rect 452542 662058 452574 662294
rect 451954 626614 452574 662058
rect 451954 626378 451986 626614
rect 452222 626378 452306 626614
rect 452542 626378 452574 626614
rect 451954 626294 452574 626378
rect 451954 626058 451986 626294
rect 452222 626058 452306 626294
rect 452542 626058 452574 626294
rect 451954 590614 452574 626058
rect 451954 590378 451986 590614
rect 452222 590378 452306 590614
rect 452542 590378 452574 590614
rect 451954 590294 452574 590378
rect 451954 590058 451986 590294
rect 452222 590058 452306 590294
rect 452542 590058 452574 590294
rect 451954 554614 452574 590058
rect 451954 554378 451986 554614
rect 452222 554378 452306 554614
rect 452542 554378 452574 554614
rect 451954 554294 452574 554378
rect 451954 554058 451986 554294
rect 452222 554058 452306 554294
rect 452542 554058 452574 554294
rect 451954 518614 452574 554058
rect 451954 518378 451986 518614
rect 452222 518378 452306 518614
rect 452542 518378 452574 518614
rect 451954 518294 452574 518378
rect 451954 518058 451986 518294
rect 452222 518058 452306 518294
rect 452542 518058 452574 518294
rect 451954 482614 452574 518058
rect 451954 482378 451986 482614
rect 452222 482378 452306 482614
rect 452542 482378 452574 482614
rect 451954 482294 452574 482378
rect 451954 482058 451986 482294
rect 452222 482058 452306 482294
rect 452542 482058 452574 482294
rect 451954 446614 452574 482058
rect 451954 446378 451986 446614
rect 452222 446378 452306 446614
rect 452542 446378 452574 446614
rect 451954 446294 452574 446378
rect 451954 446058 451986 446294
rect 452222 446058 452306 446294
rect 452542 446058 452574 446294
rect 451954 410614 452574 446058
rect 451954 410378 451986 410614
rect 452222 410378 452306 410614
rect 452542 410378 452574 410614
rect 451954 410294 452574 410378
rect 451954 410058 451986 410294
rect 452222 410058 452306 410294
rect 452542 410058 452574 410294
rect 451954 374614 452574 410058
rect 451954 374378 451986 374614
rect 452222 374378 452306 374614
rect 452542 374378 452574 374614
rect 451954 374294 452574 374378
rect 451954 374058 451986 374294
rect 452222 374058 452306 374294
rect 452542 374058 452574 374294
rect 451954 338614 452574 374058
rect 451954 338378 451986 338614
rect 452222 338378 452306 338614
rect 452542 338378 452574 338614
rect 451954 338294 452574 338378
rect 451954 338058 451986 338294
rect 452222 338058 452306 338294
rect 452542 338058 452574 338294
rect 451954 302614 452574 338058
rect 451954 302378 451986 302614
rect 452222 302378 452306 302614
rect 452542 302378 452574 302614
rect 451954 302294 452574 302378
rect 451954 302058 451986 302294
rect 452222 302058 452306 302294
rect 452542 302058 452574 302294
rect 451954 266614 452574 302058
rect 451954 266378 451986 266614
rect 452222 266378 452306 266614
rect 452542 266378 452574 266614
rect 451954 266294 452574 266378
rect 451954 266058 451986 266294
rect 452222 266058 452306 266294
rect 452542 266058 452574 266294
rect 451954 230614 452574 266058
rect 451954 230378 451986 230614
rect 452222 230378 452306 230614
rect 452542 230378 452574 230614
rect 451954 230294 452574 230378
rect 451954 230058 451986 230294
rect 452222 230058 452306 230294
rect 452542 230058 452574 230294
rect 451954 194614 452574 230058
rect 451954 194378 451986 194614
rect 452222 194378 452306 194614
rect 452542 194378 452574 194614
rect 451954 194294 452574 194378
rect 451954 194058 451986 194294
rect 452222 194058 452306 194294
rect 452542 194058 452574 194294
rect 451954 158614 452574 194058
rect 451954 158378 451986 158614
rect 452222 158378 452306 158614
rect 452542 158378 452574 158614
rect 451954 158294 452574 158378
rect 451954 158058 451986 158294
rect 452222 158058 452306 158294
rect 452542 158058 452574 158294
rect 451954 122614 452574 158058
rect 451954 122378 451986 122614
rect 452222 122378 452306 122614
rect 452542 122378 452574 122614
rect 451954 122294 452574 122378
rect 451954 122058 451986 122294
rect 452222 122058 452306 122294
rect 452542 122058 452574 122294
rect 451954 86614 452574 122058
rect 451954 86378 451986 86614
rect 452222 86378 452306 86614
rect 452542 86378 452574 86614
rect 451954 86294 452574 86378
rect 451954 86058 451986 86294
rect 452222 86058 452306 86294
rect 452542 86058 452574 86294
rect 451954 50614 452574 86058
rect 451954 50378 451986 50614
rect 452222 50378 452306 50614
rect 452542 50378 452574 50614
rect 451954 50294 452574 50378
rect 451954 50058 451986 50294
rect 452222 50058 452306 50294
rect 452542 50058 452574 50294
rect 451954 14614 452574 50058
rect 451954 14378 451986 14614
rect 452222 14378 452306 14614
rect 452542 14378 452574 14614
rect 451954 14294 452574 14378
rect 451954 14058 451986 14294
rect 452222 14058 452306 14294
rect 452542 14058 452574 14294
rect 448234 -4422 448266 -4186
rect 448502 -4422 448586 -4186
rect 448822 -4422 448854 -4186
rect 448234 -4506 448854 -4422
rect 448234 -4742 448266 -4506
rect 448502 -4742 448586 -4506
rect 448822 -4742 448854 -4506
rect 448234 -5734 448854 -4742
rect 441954 -7302 441986 -7066
rect 442222 -7302 442306 -7066
rect 442542 -7302 442574 -7066
rect 441954 -7386 442574 -7302
rect 441954 -7622 441986 -7386
rect 442222 -7622 442306 -7386
rect 442542 -7622 442574 -7386
rect 441954 -7654 442574 -7622
rect 451954 -6106 452574 14058
rect 454514 707718 455134 707750
rect 454514 707482 454546 707718
rect 454782 707482 454866 707718
rect 455102 707482 455134 707718
rect 454514 707398 455134 707482
rect 454514 707162 454546 707398
rect 454782 707162 454866 707398
rect 455102 707162 455134 707398
rect 454514 673174 455134 707162
rect 454514 672938 454546 673174
rect 454782 672938 454866 673174
rect 455102 672938 455134 673174
rect 454514 672854 455134 672938
rect 454514 672618 454546 672854
rect 454782 672618 454866 672854
rect 455102 672618 455134 672854
rect 454514 637174 455134 672618
rect 454514 636938 454546 637174
rect 454782 636938 454866 637174
rect 455102 636938 455134 637174
rect 454514 636854 455134 636938
rect 454514 636618 454546 636854
rect 454782 636618 454866 636854
rect 455102 636618 455134 636854
rect 454514 601174 455134 636618
rect 454514 600938 454546 601174
rect 454782 600938 454866 601174
rect 455102 600938 455134 601174
rect 454514 600854 455134 600938
rect 454514 600618 454546 600854
rect 454782 600618 454866 600854
rect 455102 600618 455134 600854
rect 454514 565174 455134 600618
rect 454514 564938 454546 565174
rect 454782 564938 454866 565174
rect 455102 564938 455134 565174
rect 454514 564854 455134 564938
rect 454514 564618 454546 564854
rect 454782 564618 454866 564854
rect 455102 564618 455134 564854
rect 454514 529174 455134 564618
rect 454514 528938 454546 529174
rect 454782 528938 454866 529174
rect 455102 528938 455134 529174
rect 454514 528854 455134 528938
rect 454514 528618 454546 528854
rect 454782 528618 454866 528854
rect 455102 528618 455134 528854
rect 454514 493174 455134 528618
rect 454514 492938 454546 493174
rect 454782 492938 454866 493174
rect 455102 492938 455134 493174
rect 454514 492854 455134 492938
rect 454514 492618 454546 492854
rect 454782 492618 454866 492854
rect 455102 492618 455134 492854
rect 454514 457174 455134 492618
rect 454514 456938 454546 457174
rect 454782 456938 454866 457174
rect 455102 456938 455134 457174
rect 454514 456854 455134 456938
rect 454514 456618 454546 456854
rect 454782 456618 454866 456854
rect 455102 456618 455134 456854
rect 454514 421174 455134 456618
rect 454514 420938 454546 421174
rect 454782 420938 454866 421174
rect 455102 420938 455134 421174
rect 454514 420854 455134 420938
rect 454514 420618 454546 420854
rect 454782 420618 454866 420854
rect 455102 420618 455134 420854
rect 454514 385174 455134 420618
rect 454514 384938 454546 385174
rect 454782 384938 454866 385174
rect 455102 384938 455134 385174
rect 454514 384854 455134 384938
rect 454514 384618 454546 384854
rect 454782 384618 454866 384854
rect 455102 384618 455134 384854
rect 454514 349174 455134 384618
rect 454514 348938 454546 349174
rect 454782 348938 454866 349174
rect 455102 348938 455134 349174
rect 454514 348854 455134 348938
rect 454514 348618 454546 348854
rect 454782 348618 454866 348854
rect 455102 348618 455134 348854
rect 454514 313174 455134 348618
rect 454514 312938 454546 313174
rect 454782 312938 454866 313174
rect 455102 312938 455134 313174
rect 454514 312854 455134 312938
rect 454514 312618 454546 312854
rect 454782 312618 454866 312854
rect 455102 312618 455134 312854
rect 454514 277174 455134 312618
rect 454514 276938 454546 277174
rect 454782 276938 454866 277174
rect 455102 276938 455134 277174
rect 454514 276854 455134 276938
rect 454514 276618 454546 276854
rect 454782 276618 454866 276854
rect 455102 276618 455134 276854
rect 454514 241174 455134 276618
rect 454514 240938 454546 241174
rect 454782 240938 454866 241174
rect 455102 240938 455134 241174
rect 454514 240854 455134 240938
rect 454514 240618 454546 240854
rect 454782 240618 454866 240854
rect 455102 240618 455134 240854
rect 454514 205174 455134 240618
rect 454514 204938 454546 205174
rect 454782 204938 454866 205174
rect 455102 204938 455134 205174
rect 454514 204854 455134 204938
rect 454514 204618 454546 204854
rect 454782 204618 454866 204854
rect 455102 204618 455134 204854
rect 454514 169174 455134 204618
rect 454514 168938 454546 169174
rect 454782 168938 454866 169174
rect 455102 168938 455134 169174
rect 454514 168854 455134 168938
rect 454514 168618 454546 168854
rect 454782 168618 454866 168854
rect 455102 168618 455134 168854
rect 454514 133174 455134 168618
rect 454514 132938 454546 133174
rect 454782 132938 454866 133174
rect 455102 132938 455134 133174
rect 454514 132854 455134 132938
rect 454514 132618 454546 132854
rect 454782 132618 454866 132854
rect 455102 132618 455134 132854
rect 454514 97174 455134 132618
rect 454514 96938 454546 97174
rect 454782 96938 454866 97174
rect 455102 96938 455134 97174
rect 454514 96854 455134 96938
rect 454514 96618 454546 96854
rect 454782 96618 454866 96854
rect 455102 96618 455134 96854
rect 454514 61174 455134 96618
rect 454514 60938 454546 61174
rect 454782 60938 454866 61174
rect 455102 60938 455134 61174
rect 454514 60854 455134 60938
rect 454514 60618 454546 60854
rect 454782 60618 454866 60854
rect 455102 60618 455134 60854
rect 454514 25174 455134 60618
rect 454514 24938 454546 25174
rect 454782 24938 454866 25174
rect 455102 24938 455134 25174
rect 454514 24854 455134 24938
rect 454514 24618 454546 24854
rect 454782 24618 454866 24854
rect 455102 24618 455134 24854
rect 454514 -3226 455134 24618
rect 454514 -3462 454546 -3226
rect 454782 -3462 454866 -3226
rect 455102 -3462 455134 -3226
rect 454514 -3546 455134 -3462
rect 454514 -3782 454546 -3546
rect 454782 -3782 454866 -3546
rect 455102 -3782 455134 -3546
rect 454514 -3814 455134 -3782
rect 458234 676894 458854 709082
rect 458234 676658 458266 676894
rect 458502 676658 458586 676894
rect 458822 676658 458854 676894
rect 458234 676574 458854 676658
rect 458234 676338 458266 676574
rect 458502 676338 458586 676574
rect 458822 676338 458854 676574
rect 458234 640894 458854 676338
rect 458234 640658 458266 640894
rect 458502 640658 458586 640894
rect 458822 640658 458854 640894
rect 458234 640574 458854 640658
rect 458234 640338 458266 640574
rect 458502 640338 458586 640574
rect 458822 640338 458854 640574
rect 458234 604894 458854 640338
rect 458234 604658 458266 604894
rect 458502 604658 458586 604894
rect 458822 604658 458854 604894
rect 458234 604574 458854 604658
rect 458234 604338 458266 604574
rect 458502 604338 458586 604574
rect 458822 604338 458854 604574
rect 458234 568894 458854 604338
rect 458234 568658 458266 568894
rect 458502 568658 458586 568894
rect 458822 568658 458854 568894
rect 458234 568574 458854 568658
rect 458234 568338 458266 568574
rect 458502 568338 458586 568574
rect 458822 568338 458854 568574
rect 458234 532894 458854 568338
rect 458234 532658 458266 532894
rect 458502 532658 458586 532894
rect 458822 532658 458854 532894
rect 458234 532574 458854 532658
rect 458234 532338 458266 532574
rect 458502 532338 458586 532574
rect 458822 532338 458854 532574
rect 458234 496894 458854 532338
rect 458234 496658 458266 496894
rect 458502 496658 458586 496894
rect 458822 496658 458854 496894
rect 458234 496574 458854 496658
rect 458234 496338 458266 496574
rect 458502 496338 458586 496574
rect 458822 496338 458854 496574
rect 458234 460894 458854 496338
rect 458234 460658 458266 460894
rect 458502 460658 458586 460894
rect 458822 460658 458854 460894
rect 458234 460574 458854 460658
rect 458234 460338 458266 460574
rect 458502 460338 458586 460574
rect 458822 460338 458854 460574
rect 458234 424894 458854 460338
rect 458234 424658 458266 424894
rect 458502 424658 458586 424894
rect 458822 424658 458854 424894
rect 458234 424574 458854 424658
rect 458234 424338 458266 424574
rect 458502 424338 458586 424574
rect 458822 424338 458854 424574
rect 458234 388894 458854 424338
rect 458234 388658 458266 388894
rect 458502 388658 458586 388894
rect 458822 388658 458854 388894
rect 458234 388574 458854 388658
rect 458234 388338 458266 388574
rect 458502 388338 458586 388574
rect 458822 388338 458854 388574
rect 458234 352894 458854 388338
rect 458234 352658 458266 352894
rect 458502 352658 458586 352894
rect 458822 352658 458854 352894
rect 458234 352574 458854 352658
rect 458234 352338 458266 352574
rect 458502 352338 458586 352574
rect 458822 352338 458854 352574
rect 458234 316894 458854 352338
rect 458234 316658 458266 316894
rect 458502 316658 458586 316894
rect 458822 316658 458854 316894
rect 458234 316574 458854 316658
rect 458234 316338 458266 316574
rect 458502 316338 458586 316574
rect 458822 316338 458854 316574
rect 458234 280894 458854 316338
rect 458234 280658 458266 280894
rect 458502 280658 458586 280894
rect 458822 280658 458854 280894
rect 458234 280574 458854 280658
rect 458234 280338 458266 280574
rect 458502 280338 458586 280574
rect 458822 280338 458854 280574
rect 458234 244894 458854 280338
rect 458234 244658 458266 244894
rect 458502 244658 458586 244894
rect 458822 244658 458854 244894
rect 458234 244574 458854 244658
rect 458234 244338 458266 244574
rect 458502 244338 458586 244574
rect 458822 244338 458854 244574
rect 458234 208894 458854 244338
rect 458234 208658 458266 208894
rect 458502 208658 458586 208894
rect 458822 208658 458854 208894
rect 458234 208574 458854 208658
rect 458234 208338 458266 208574
rect 458502 208338 458586 208574
rect 458822 208338 458854 208574
rect 458234 172894 458854 208338
rect 458234 172658 458266 172894
rect 458502 172658 458586 172894
rect 458822 172658 458854 172894
rect 458234 172574 458854 172658
rect 458234 172338 458266 172574
rect 458502 172338 458586 172574
rect 458822 172338 458854 172574
rect 458234 136894 458854 172338
rect 458234 136658 458266 136894
rect 458502 136658 458586 136894
rect 458822 136658 458854 136894
rect 458234 136574 458854 136658
rect 458234 136338 458266 136574
rect 458502 136338 458586 136574
rect 458822 136338 458854 136574
rect 458234 100894 458854 136338
rect 458234 100658 458266 100894
rect 458502 100658 458586 100894
rect 458822 100658 458854 100894
rect 458234 100574 458854 100658
rect 458234 100338 458266 100574
rect 458502 100338 458586 100574
rect 458822 100338 458854 100574
rect 458234 64894 458854 100338
rect 458234 64658 458266 64894
rect 458502 64658 458586 64894
rect 458822 64658 458854 64894
rect 458234 64574 458854 64658
rect 458234 64338 458266 64574
rect 458502 64338 458586 64574
rect 458822 64338 458854 64574
rect 458234 28894 458854 64338
rect 458234 28658 458266 28894
rect 458502 28658 458586 28894
rect 458822 28658 458854 28894
rect 458234 28574 458854 28658
rect 458234 28338 458266 28574
rect 458502 28338 458586 28574
rect 458822 28338 458854 28574
rect 458234 -5146 458854 28338
rect 460794 704838 461414 705830
rect 460794 704602 460826 704838
rect 461062 704602 461146 704838
rect 461382 704602 461414 704838
rect 460794 704518 461414 704602
rect 460794 704282 460826 704518
rect 461062 704282 461146 704518
rect 461382 704282 461414 704518
rect 460794 687454 461414 704282
rect 460794 687218 460826 687454
rect 461062 687218 461146 687454
rect 461382 687218 461414 687454
rect 460794 687134 461414 687218
rect 460794 686898 460826 687134
rect 461062 686898 461146 687134
rect 461382 686898 461414 687134
rect 460794 651454 461414 686898
rect 460794 651218 460826 651454
rect 461062 651218 461146 651454
rect 461382 651218 461414 651454
rect 460794 651134 461414 651218
rect 460794 650898 460826 651134
rect 461062 650898 461146 651134
rect 461382 650898 461414 651134
rect 460794 615454 461414 650898
rect 460794 615218 460826 615454
rect 461062 615218 461146 615454
rect 461382 615218 461414 615454
rect 460794 615134 461414 615218
rect 460794 614898 460826 615134
rect 461062 614898 461146 615134
rect 461382 614898 461414 615134
rect 460794 579454 461414 614898
rect 460794 579218 460826 579454
rect 461062 579218 461146 579454
rect 461382 579218 461414 579454
rect 460794 579134 461414 579218
rect 460794 578898 460826 579134
rect 461062 578898 461146 579134
rect 461382 578898 461414 579134
rect 460794 543454 461414 578898
rect 460794 543218 460826 543454
rect 461062 543218 461146 543454
rect 461382 543218 461414 543454
rect 460794 543134 461414 543218
rect 460794 542898 460826 543134
rect 461062 542898 461146 543134
rect 461382 542898 461414 543134
rect 460794 507454 461414 542898
rect 460794 507218 460826 507454
rect 461062 507218 461146 507454
rect 461382 507218 461414 507454
rect 460794 507134 461414 507218
rect 460794 506898 460826 507134
rect 461062 506898 461146 507134
rect 461382 506898 461414 507134
rect 460794 471454 461414 506898
rect 460794 471218 460826 471454
rect 461062 471218 461146 471454
rect 461382 471218 461414 471454
rect 460794 471134 461414 471218
rect 460794 470898 460826 471134
rect 461062 470898 461146 471134
rect 461382 470898 461414 471134
rect 460794 435454 461414 470898
rect 460794 435218 460826 435454
rect 461062 435218 461146 435454
rect 461382 435218 461414 435454
rect 460794 435134 461414 435218
rect 460794 434898 460826 435134
rect 461062 434898 461146 435134
rect 461382 434898 461414 435134
rect 460794 399454 461414 434898
rect 460794 399218 460826 399454
rect 461062 399218 461146 399454
rect 461382 399218 461414 399454
rect 460794 399134 461414 399218
rect 460794 398898 460826 399134
rect 461062 398898 461146 399134
rect 461382 398898 461414 399134
rect 460794 363454 461414 398898
rect 460794 363218 460826 363454
rect 461062 363218 461146 363454
rect 461382 363218 461414 363454
rect 460794 363134 461414 363218
rect 460794 362898 460826 363134
rect 461062 362898 461146 363134
rect 461382 362898 461414 363134
rect 460794 327454 461414 362898
rect 460794 327218 460826 327454
rect 461062 327218 461146 327454
rect 461382 327218 461414 327454
rect 460794 327134 461414 327218
rect 460794 326898 460826 327134
rect 461062 326898 461146 327134
rect 461382 326898 461414 327134
rect 460794 291454 461414 326898
rect 460794 291218 460826 291454
rect 461062 291218 461146 291454
rect 461382 291218 461414 291454
rect 460794 291134 461414 291218
rect 460794 290898 460826 291134
rect 461062 290898 461146 291134
rect 461382 290898 461414 291134
rect 460794 255454 461414 290898
rect 460794 255218 460826 255454
rect 461062 255218 461146 255454
rect 461382 255218 461414 255454
rect 460794 255134 461414 255218
rect 460794 254898 460826 255134
rect 461062 254898 461146 255134
rect 461382 254898 461414 255134
rect 460794 219454 461414 254898
rect 460794 219218 460826 219454
rect 461062 219218 461146 219454
rect 461382 219218 461414 219454
rect 460794 219134 461414 219218
rect 460794 218898 460826 219134
rect 461062 218898 461146 219134
rect 461382 218898 461414 219134
rect 460794 183454 461414 218898
rect 460794 183218 460826 183454
rect 461062 183218 461146 183454
rect 461382 183218 461414 183454
rect 460794 183134 461414 183218
rect 460794 182898 460826 183134
rect 461062 182898 461146 183134
rect 461382 182898 461414 183134
rect 460794 147454 461414 182898
rect 460794 147218 460826 147454
rect 461062 147218 461146 147454
rect 461382 147218 461414 147454
rect 460794 147134 461414 147218
rect 460794 146898 460826 147134
rect 461062 146898 461146 147134
rect 461382 146898 461414 147134
rect 460794 111454 461414 146898
rect 460794 111218 460826 111454
rect 461062 111218 461146 111454
rect 461382 111218 461414 111454
rect 460794 111134 461414 111218
rect 460794 110898 460826 111134
rect 461062 110898 461146 111134
rect 461382 110898 461414 111134
rect 460794 75454 461414 110898
rect 460794 75218 460826 75454
rect 461062 75218 461146 75454
rect 461382 75218 461414 75454
rect 460794 75134 461414 75218
rect 460794 74898 460826 75134
rect 461062 74898 461146 75134
rect 461382 74898 461414 75134
rect 460794 39454 461414 74898
rect 460794 39218 460826 39454
rect 461062 39218 461146 39454
rect 461382 39218 461414 39454
rect 460794 39134 461414 39218
rect 460794 38898 460826 39134
rect 461062 38898 461146 39134
rect 461382 38898 461414 39134
rect 460794 3454 461414 38898
rect 460794 3218 460826 3454
rect 461062 3218 461146 3454
rect 461382 3218 461414 3454
rect 460794 3134 461414 3218
rect 460794 2898 460826 3134
rect 461062 2898 461146 3134
rect 461382 2898 461414 3134
rect 460794 -346 461414 2898
rect 460794 -582 460826 -346
rect 461062 -582 461146 -346
rect 461382 -582 461414 -346
rect 460794 -666 461414 -582
rect 460794 -902 460826 -666
rect 461062 -902 461146 -666
rect 461382 -902 461414 -666
rect 460794 -1894 461414 -902
rect 461954 680614 462574 711002
rect 471954 710598 472574 711590
rect 471954 710362 471986 710598
rect 472222 710362 472306 710598
rect 472542 710362 472574 710598
rect 471954 710278 472574 710362
rect 471954 710042 471986 710278
rect 472222 710042 472306 710278
rect 472542 710042 472574 710278
rect 468234 708678 468854 709670
rect 468234 708442 468266 708678
rect 468502 708442 468586 708678
rect 468822 708442 468854 708678
rect 468234 708358 468854 708442
rect 468234 708122 468266 708358
rect 468502 708122 468586 708358
rect 468822 708122 468854 708358
rect 461954 680378 461986 680614
rect 462222 680378 462306 680614
rect 462542 680378 462574 680614
rect 461954 680294 462574 680378
rect 461954 680058 461986 680294
rect 462222 680058 462306 680294
rect 462542 680058 462574 680294
rect 461954 644614 462574 680058
rect 461954 644378 461986 644614
rect 462222 644378 462306 644614
rect 462542 644378 462574 644614
rect 461954 644294 462574 644378
rect 461954 644058 461986 644294
rect 462222 644058 462306 644294
rect 462542 644058 462574 644294
rect 461954 608614 462574 644058
rect 461954 608378 461986 608614
rect 462222 608378 462306 608614
rect 462542 608378 462574 608614
rect 461954 608294 462574 608378
rect 461954 608058 461986 608294
rect 462222 608058 462306 608294
rect 462542 608058 462574 608294
rect 461954 572614 462574 608058
rect 461954 572378 461986 572614
rect 462222 572378 462306 572614
rect 462542 572378 462574 572614
rect 461954 572294 462574 572378
rect 461954 572058 461986 572294
rect 462222 572058 462306 572294
rect 462542 572058 462574 572294
rect 461954 536614 462574 572058
rect 461954 536378 461986 536614
rect 462222 536378 462306 536614
rect 462542 536378 462574 536614
rect 461954 536294 462574 536378
rect 461954 536058 461986 536294
rect 462222 536058 462306 536294
rect 462542 536058 462574 536294
rect 461954 500614 462574 536058
rect 461954 500378 461986 500614
rect 462222 500378 462306 500614
rect 462542 500378 462574 500614
rect 461954 500294 462574 500378
rect 461954 500058 461986 500294
rect 462222 500058 462306 500294
rect 462542 500058 462574 500294
rect 461954 464614 462574 500058
rect 461954 464378 461986 464614
rect 462222 464378 462306 464614
rect 462542 464378 462574 464614
rect 461954 464294 462574 464378
rect 461954 464058 461986 464294
rect 462222 464058 462306 464294
rect 462542 464058 462574 464294
rect 461954 428614 462574 464058
rect 461954 428378 461986 428614
rect 462222 428378 462306 428614
rect 462542 428378 462574 428614
rect 461954 428294 462574 428378
rect 461954 428058 461986 428294
rect 462222 428058 462306 428294
rect 462542 428058 462574 428294
rect 461954 392614 462574 428058
rect 461954 392378 461986 392614
rect 462222 392378 462306 392614
rect 462542 392378 462574 392614
rect 461954 392294 462574 392378
rect 461954 392058 461986 392294
rect 462222 392058 462306 392294
rect 462542 392058 462574 392294
rect 461954 356614 462574 392058
rect 461954 356378 461986 356614
rect 462222 356378 462306 356614
rect 462542 356378 462574 356614
rect 461954 356294 462574 356378
rect 461954 356058 461986 356294
rect 462222 356058 462306 356294
rect 462542 356058 462574 356294
rect 461954 320614 462574 356058
rect 461954 320378 461986 320614
rect 462222 320378 462306 320614
rect 462542 320378 462574 320614
rect 461954 320294 462574 320378
rect 461954 320058 461986 320294
rect 462222 320058 462306 320294
rect 462542 320058 462574 320294
rect 461954 284614 462574 320058
rect 461954 284378 461986 284614
rect 462222 284378 462306 284614
rect 462542 284378 462574 284614
rect 461954 284294 462574 284378
rect 461954 284058 461986 284294
rect 462222 284058 462306 284294
rect 462542 284058 462574 284294
rect 461954 248614 462574 284058
rect 461954 248378 461986 248614
rect 462222 248378 462306 248614
rect 462542 248378 462574 248614
rect 461954 248294 462574 248378
rect 461954 248058 461986 248294
rect 462222 248058 462306 248294
rect 462542 248058 462574 248294
rect 461954 212614 462574 248058
rect 461954 212378 461986 212614
rect 462222 212378 462306 212614
rect 462542 212378 462574 212614
rect 461954 212294 462574 212378
rect 461954 212058 461986 212294
rect 462222 212058 462306 212294
rect 462542 212058 462574 212294
rect 461954 176614 462574 212058
rect 461954 176378 461986 176614
rect 462222 176378 462306 176614
rect 462542 176378 462574 176614
rect 461954 176294 462574 176378
rect 461954 176058 461986 176294
rect 462222 176058 462306 176294
rect 462542 176058 462574 176294
rect 461954 140614 462574 176058
rect 461954 140378 461986 140614
rect 462222 140378 462306 140614
rect 462542 140378 462574 140614
rect 461954 140294 462574 140378
rect 461954 140058 461986 140294
rect 462222 140058 462306 140294
rect 462542 140058 462574 140294
rect 461954 104614 462574 140058
rect 461954 104378 461986 104614
rect 462222 104378 462306 104614
rect 462542 104378 462574 104614
rect 461954 104294 462574 104378
rect 461954 104058 461986 104294
rect 462222 104058 462306 104294
rect 462542 104058 462574 104294
rect 461954 68614 462574 104058
rect 461954 68378 461986 68614
rect 462222 68378 462306 68614
rect 462542 68378 462574 68614
rect 461954 68294 462574 68378
rect 461954 68058 461986 68294
rect 462222 68058 462306 68294
rect 462542 68058 462574 68294
rect 461954 32614 462574 68058
rect 461954 32378 461986 32614
rect 462222 32378 462306 32614
rect 462542 32378 462574 32614
rect 461954 32294 462574 32378
rect 461954 32058 461986 32294
rect 462222 32058 462306 32294
rect 462542 32058 462574 32294
rect 458234 -5382 458266 -5146
rect 458502 -5382 458586 -5146
rect 458822 -5382 458854 -5146
rect 458234 -5466 458854 -5382
rect 458234 -5702 458266 -5466
rect 458502 -5702 458586 -5466
rect 458822 -5702 458854 -5466
rect 458234 -5734 458854 -5702
rect 451954 -6342 451986 -6106
rect 452222 -6342 452306 -6106
rect 452542 -6342 452574 -6106
rect 451954 -6426 452574 -6342
rect 451954 -6662 451986 -6426
rect 452222 -6662 452306 -6426
rect 452542 -6662 452574 -6426
rect 451954 -7654 452574 -6662
rect 461954 -7066 462574 32058
rect 464514 706758 465134 707750
rect 464514 706522 464546 706758
rect 464782 706522 464866 706758
rect 465102 706522 465134 706758
rect 464514 706438 465134 706522
rect 464514 706202 464546 706438
rect 464782 706202 464866 706438
rect 465102 706202 465134 706438
rect 464514 691174 465134 706202
rect 464514 690938 464546 691174
rect 464782 690938 464866 691174
rect 465102 690938 465134 691174
rect 464514 690854 465134 690938
rect 464514 690618 464546 690854
rect 464782 690618 464866 690854
rect 465102 690618 465134 690854
rect 464514 655174 465134 690618
rect 464514 654938 464546 655174
rect 464782 654938 464866 655174
rect 465102 654938 465134 655174
rect 464514 654854 465134 654938
rect 464514 654618 464546 654854
rect 464782 654618 464866 654854
rect 465102 654618 465134 654854
rect 464514 619174 465134 654618
rect 464514 618938 464546 619174
rect 464782 618938 464866 619174
rect 465102 618938 465134 619174
rect 464514 618854 465134 618938
rect 464514 618618 464546 618854
rect 464782 618618 464866 618854
rect 465102 618618 465134 618854
rect 464514 583174 465134 618618
rect 464514 582938 464546 583174
rect 464782 582938 464866 583174
rect 465102 582938 465134 583174
rect 464514 582854 465134 582938
rect 464514 582618 464546 582854
rect 464782 582618 464866 582854
rect 465102 582618 465134 582854
rect 464514 547174 465134 582618
rect 464514 546938 464546 547174
rect 464782 546938 464866 547174
rect 465102 546938 465134 547174
rect 464514 546854 465134 546938
rect 464514 546618 464546 546854
rect 464782 546618 464866 546854
rect 465102 546618 465134 546854
rect 464514 511174 465134 546618
rect 464514 510938 464546 511174
rect 464782 510938 464866 511174
rect 465102 510938 465134 511174
rect 464514 510854 465134 510938
rect 464514 510618 464546 510854
rect 464782 510618 464866 510854
rect 465102 510618 465134 510854
rect 464514 475174 465134 510618
rect 464514 474938 464546 475174
rect 464782 474938 464866 475174
rect 465102 474938 465134 475174
rect 464514 474854 465134 474938
rect 464514 474618 464546 474854
rect 464782 474618 464866 474854
rect 465102 474618 465134 474854
rect 464514 439174 465134 474618
rect 464514 438938 464546 439174
rect 464782 438938 464866 439174
rect 465102 438938 465134 439174
rect 464514 438854 465134 438938
rect 464514 438618 464546 438854
rect 464782 438618 464866 438854
rect 465102 438618 465134 438854
rect 464514 403174 465134 438618
rect 464514 402938 464546 403174
rect 464782 402938 464866 403174
rect 465102 402938 465134 403174
rect 464514 402854 465134 402938
rect 464514 402618 464546 402854
rect 464782 402618 464866 402854
rect 465102 402618 465134 402854
rect 464514 367174 465134 402618
rect 464514 366938 464546 367174
rect 464782 366938 464866 367174
rect 465102 366938 465134 367174
rect 464514 366854 465134 366938
rect 464514 366618 464546 366854
rect 464782 366618 464866 366854
rect 465102 366618 465134 366854
rect 464514 331174 465134 366618
rect 464514 330938 464546 331174
rect 464782 330938 464866 331174
rect 465102 330938 465134 331174
rect 464514 330854 465134 330938
rect 464514 330618 464546 330854
rect 464782 330618 464866 330854
rect 465102 330618 465134 330854
rect 464514 295174 465134 330618
rect 464514 294938 464546 295174
rect 464782 294938 464866 295174
rect 465102 294938 465134 295174
rect 464514 294854 465134 294938
rect 464514 294618 464546 294854
rect 464782 294618 464866 294854
rect 465102 294618 465134 294854
rect 464514 259174 465134 294618
rect 464514 258938 464546 259174
rect 464782 258938 464866 259174
rect 465102 258938 465134 259174
rect 464514 258854 465134 258938
rect 464514 258618 464546 258854
rect 464782 258618 464866 258854
rect 465102 258618 465134 258854
rect 464514 223174 465134 258618
rect 464514 222938 464546 223174
rect 464782 222938 464866 223174
rect 465102 222938 465134 223174
rect 464514 222854 465134 222938
rect 464514 222618 464546 222854
rect 464782 222618 464866 222854
rect 465102 222618 465134 222854
rect 464514 187174 465134 222618
rect 464514 186938 464546 187174
rect 464782 186938 464866 187174
rect 465102 186938 465134 187174
rect 464514 186854 465134 186938
rect 464514 186618 464546 186854
rect 464782 186618 464866 186854
rect 465102 186618 465134 186854
rect 464514 151174 465134 186618
rect 464514 150938 464546 151174
rect 464782 150938 464866 151174
rect 465102 150938 465134 151174
rect 464514 150854 465134 150938
rect 464514 150618 464546 150854
rect 464782 150618 464866 150854
rect 465102 150618 465134 150854
rect 464514 115174 465134 150618
rect 464514 114938 464546 115174
rect 464782 114938 464866 115174
rect 465102 114938 465134 115174
rect 464514 114854 465134 114938
rect 464514 114618 464546 114854
rect 464782 114618 464866 114854
rect 465102 114618 465134 114854
rect 464514 79174 465134 114618
rect 464514 78938 464546 79174
rect 464782 78938 464866 79174
rect 465102 78938 465134 79174
rect 464514 78854 465134 78938
rect 464514 78618 464546 78854
rect 464782 78618 464866 78854
rect 465102 78618 465134 78854
rect 464514 43174 465134 78618
rect 464514 42938 464546 43174
rect 464782 42938 464866 43174
rect 465102 42938 465134 43174
rect 464514 42854 465134 42938
rect 464514 42618 464546 42854
rect 464782 42618 464866 42854
rect 465102 42618 465134 42854
rect 464514 7174 465134 42618
rect 464514 6938 464546 7174
rect 464782 6938 464866 7174
rect 465102 6938 465134 7174
rect 464514 6854 465134 6938
rect 464514 6618 464546 6854
rect 464782 6618 464866 6854
rect 465102 6618 465134 6854
rect 464514 -2266 465134 6618
rect 464514 -2502 464546 -2266
rect 464782 -2502 464866 -2266
rect 465102 -2502 465134 -2266
rect 464514 -2586 465134 -2502
rect 464514 -2822 464546 -2586
rect 464782 -2822 464866 -2586
rect 465102 -2822 465134 -2586
rect 464514 -3814 465134 -2822
rect 468234 694894 468854 708122
rect 468234 694658 468266 694894
rect 468502 694658 468586 694894
rect 468822 694658 468854 694894
rect 468234 694574 468854 694658
rect 468234 694338 468266 694574
rect 468502 694338 468586 694574
rect 468822 694338 468854 694574
rect 468234 658894 468854 694338
rect 468234 658658 468266 658894
rect 468502 658658 468586 658894
rect 468822 658658 468854 658894
rect 468234 658574 468854 658658
rect 468234 658338 468266 658574
rect 468502 658338 468586 658574
rect 468822 658338 468854 658574
rect 468234 622894 468854 658338
rect 468234 622658 468266 622894
rect 468502 622658 468586 622894
rect 468822 622658 468854 622894
rect 468234 622574 468854 622658
rect 468234 622338 468266 622574
rect 468502 622338 468586 622574
rect 468822 622338 468854 622574
rect 468234 586894 468854 622338
rect 468234 586658 468266 586894
rect 468502 586658 468586 586894
rect 468822 586658 468854 586894
rect 468234 586574 468854 586658
rect 468234 586338 468266 586574
rect 468502 586338 468586 586574
rect 468822 586338 468854 586574
rect 468234 550894 468854 586338
rect 468234 550658 468266 550894
rect 468502 550658 468586 550894
rect 468822 550658 468854 550894
rect 468234 550574 468854 550658
rect 468234 550338 468266 550574
rect 468502 550338 468586 550574
rect 468822 550338 468854 550574
rect 468234 514894 468854 550338
rect 468234 514658 468266 514894
rect 468502 514658 468586 514894
rect 468822 514658 468854 514894
rect 468234 514574 468854 514658
rect 468234 514338 468266 514574
rect 468502 514338 468586 514574
rect 468822 514338 468854 514574
rect 468234 478894 468854 514338
rect 468234 478658 468266 478894
rect 468502 478658 468586 478894
rect 468822 478658 468854 478894
rect 468234 478574 468854 478658
rect 468234 478338 468266 478574
rect 468502 478338 468586 478574
rect 468822 478338 468854 478574
rect 468234 442894 468854 478338
rect 468234 442658 468266 442894
rect 468502 442658 468586 442894
rect 468822 442658 468854 442894
rect 468234 442574 468854 442658
rect 468234 442338 468266 442574
rect 468502 442338 468586 442574
rect 468822 442338 468854 442574
rect 468234 406894 468854 442338
rect 468234 406658 468266 406894
rect 468502 406658 468586 406894
rect 468822 406658 468854 406894
rect 468234 406574 468854 406658
rect 468234 406338 468266 406574
rect 468502 406338 468586 406574
rect 468822 406338 468854 406574
rect 468234 370894 468854 406338
rect 468234 370658 468266 370894
rect 468502 370658 468586 370894
rect 468822 370658 468854 370894
rect 468234 370574 468854 370658
rect 468234 370338 468266 370574
rect 468502 370338 468586 370574
rect 468822 370338 468854 370574
rect 468234 334894 468854 370338
rect 468234 334658 468266 334894
rect 468502 334658 468586 334894
rect 468822 334658 468854 334894
rect 468234 334574 468854 334658
rect 468234 334338 468266 334574
rect 468502 334338 468586 334574
rect 468822 334338 468854 334574
rect 468234 298894 468854 334338
rect 468234 298658 468266 298894
rect 468502 298658 468586 298894
rect 468822 298658 468854 298894
rect 468234 298574 468854 298658
rect 468234 298338 468266 298574
rect 468502 298338 468586 298574
rect 468822 298338 468854 298574
rect 468234 262894 468854 298338
rect 468234 262658 468266 262894
rect 468502 262658 468586 262894
rect 468822 262658 468854 262894
rect 468234 262574 468854 262658
rect 468234 262338 468266 262574
rect 468502 262338 468586 262574
rect 468822 262338 468854 262574
rect 468234 226894 468854 262338
rect 468234 226658 468266 226894
rect 468502 226658 468586 226894
rect 468822 226658 468854 226894
rect 468234 226574 468854 226658
rect 468234 226338 468266 226574
rect 468502 226338 468586 226574
rect 468822 226338 468854 226574
rect 468234 190894 468854 226338
rect 468234 190658 468266 190894
rect 468502 190658 468586 190894
rect 468822 190658 468854 190894
rect 468234 190574 468854 190658
rect 468234 190338 468266 190574
rect 468502 190338 468586 190574
rect 468822 190338 468854 190574
rect 468234 154894 468854 190338
rect 468234 154658 468266 154894
rect 468502 154658 468586 154894
rect 468822 154658 468854 154894
rect 468234 154574 468854 154658
rect 468234 154338 468266 154574
rect 468502 154338 468586 154574
rect 468822 154338 468854 154574
rect 468234 118894 468854 154338
rect 468234 118658 468266 118894
rect 468502 118658 468586 118894
rect 468822 118658 468854 118894
rect 468234 118574 468854 118658
rect 468234 118338 468266 118574
rect 468502 118338 468586 118574
rect 468822 118338 468854 118574
rect 468234 82894 468854 118338
rect 468234 82658 468266 82894
rect 468502 82658 468586 82894
rect 468822 82658 468854 82894
rect 468234 82574 468854 82658
rect 468234 82338 468266 82574
rect 468502 82338 468586 82574
rect 468822 82338 468854 82574
rect 468234 46894 468854 82338
rect 468234 46658 468266 46894
rect 468502 46658 468586 46894
rect 468822 46658 468854 46894
rect 468234 46574 468854 46658
rect 468234 46338 468266 46574
rect 468502 46338 468586 46574
rect 468822 46338 468854 46574
rect 468234 10894 468854 46338
rect 468234 10658 468266 10894
rect 468502 10658 468586 10894
rect 468822 10658 468854 10894
rect 468234 10574 468854 10658
rect 468234 10338 468266 10574
rect 468502 10338 468586 10574
rect 468822 10338 468854 10574
rect 468234 -4186 468854 10338
rect 470794 705798 471414 705830
rect 470794 705562 470826 705798
rect 471062 705562 471146 705798
rect 471382 705562 471414 705798
rect 470794 705478 471414 705562
rect 470794 705242 470826 705478
rect 471062 705242 471146 705478
rect 471382 705242 471414 705478
rect 470794 669454 471414 705242
rect 470794 669218 470826 669454
rect 471062 669218 471146 669454
rect 471382 669218 471414 669454
rect 470794 669134 471414 669218
rect 470794 668898 470826 669134
rect 471062 668898 471146 669134
rect 471382 668898 471414 669134
rect 470794 633454 471414 668898
rect 470794 633218 470826 633454
rect 471062 633218 471146 633454
rect 471382 633218 471414 633454
rect 470794 633134 471414 633218
rect 470794 632898 470826 633134
rect 471062 632898 471146 633134
rect 471382 632898 471414 633134
rect 470794 597454 471414 632898
rect 470794 597218 470826 597454
rect 471062 597218 471146 597454
rect 471382 597218 471414 597454
rect 470794 597134 471414 597218
rect 470794 596898 470826 597134
rect 471062 596898 471146 597134
rect 471382 596898 471414 597134
rect 470794 561454 471414 596898
rect 470794 561218 470826 561454
rect 471062 561218 471146 561454
rect 471382 561218 471414 561454
rect 470794 561134 471414 561218
rect 470794 560898 470826 561134
rect 471062 560898 471146 561134
rect 471382 560898 471414 561134
rect 470794 525454 471414 560898
rect 470794 525218 470826 525454
rect 471062 525218 471146 525454
rect 471382 525218 471414 525454
rect 470794 525134 471414 525218
rect 470794 524898 470826 525134
rect 471062 524898 471146 525134
rect 471382 524898 471414 525134
rect 470794 489454 471414 524898
rect 470794 489218 470826 489454
rect 471062 489218 471146 489454
rect 471382 489218 471414 489454
rect 470794 489134 471414 489218
rect 470794 488898 470826 489134
rect 471062 488898 471146 489134
rect 471382 488898 471414 489134
rect 470794 453454 471414 488898
rect 470794 453218 470826 453454
rect 471062 453218 471146 453454
rect 471382 453218 471414 453454
rect 470794 453134 471414 453218
rect 470794 452898 470826 453134
rect 471062 452898 471146 453134
rect 471382 452898 471414 453134
rect 470794 417454 471414 452898
rect 470794 417218 470826 417454
rect 471062 417218 471146 417454
rect 471382 417218 471414 417454
rect 470794 417134 471414 417218
rect 470794 416898 470826 417134
rect 471062 416898 471146 417134
rect 471382 416898 471414 417134
rect 470794 381454 471414 416898
rect 470794 381218 470826 381454
rect 471062 381218 471146 381454
rect 471382 381218 471414 381454
rect 470794 381134 471414 381218
rect 470794 380898 470826 381134
rect 471062 380898 471146 381134
rect 471382 380898 471414 381134
rect 470794 345454 471414 380898
rect 470794 345218 470826 345454
rect 471062 345218 471146 345454
rect 471382 345218 471414 345454
rect 470794 345134 471414 345218
rect 470794 344898 470826 345134
rect 471062 344898 471146 345134
rect 471382 344898 471414 345134
rect 470794 309454 471414 344898
rect 470794 309218 470826 309454
rect 471062 309218 471146 309454
rect 471382 309218 471414 309454
rect 470794 309134 471414 309218
rect 470794 308898 470826 309134
rect 471062 308898 471146 309134
rect 471382 308898 471414 309134
rect 470794 273454 471414 308898
rect 470794 273218 470826 273454
rect 471062 273218 471146 273454
rect 471382 273218 471414 273454
rect 470794 273134 471414 273218
rect 470794 272898 470826 273134
rect 471062 272898 471146 273134
rect 471382 272898 471414 273134
rect 470794 237454 471414 272898
rect 470794 237218 470826 237454
rect 471062 237218 471146 237454
rect 471382 237218 471414 237454
rect 470794 237134 471414 237218
rect 470794 236898 470826 237134
rect 471062 236898 471146 237134
rect 471382 236898 471414 237134
rect 470794 201454 471414 236898
rect 470794 201218 470826 201454
rect 471062 201218 471146 201454
rect 471382 201218 471414 201454
rect 470794 201134 471414 201218
rect 470794 200898 470826 201134
rect 471062 200898 471146 201134
rect 471382 200898 471414 201134
rect 470794 165454 471414 200898
rect 470794 165218 470826 165454
rect 471062 165218 471146 165454
rect 471382 165218 471414 165454
rect 470794 165134 471414 165218
rect 470794 164898 470826 165134
rect 471062 164898 471146 165134
rect 471382 164898 471414 165134
rect 470794 129454 471414 164898
rect 470794 129218 470826 129454
rect 471062 129218 471146 129454
rect 471382 129218 471414 129454
rect 470794 129134 471414 129218
rect 470794 128898 470826 129134
rect 471062 128898 471146 129134
rect 471382 128898 471414 129134
rect 470794 93454 471414 128898
rect 470794 93218 470826 93454
rect 471062 93218 471146 93454
rect 471382 93218 471414 93454
rect 470794 93134 471414 93218
rect 470794 92898 470826 93134
rect 471062 92898 471146 93134
rect 471382 92898 471414 93134
rect 470794 57454 471414 92898
rect 470794 57218 470826 57454
rect 471062 57218 471146 57454
rect 471382 57218 471414 57454
rect 470794 57134 471414 57218
rect 470794 56898 470826 57134
rect 471062 56898 471146 57134
rect 471382 56898 471414 57134
rect 470794 21454 471414 56898
rect 470794 21218 470826 21454
rect 471062 21218 471146 21454
rect 471382 21218 471414 21454
rect 470794 21134 471414 21218
rect 470794 20898 470826 21134
rect 471062 20898 471146 21134
rect 471382 20898 471414 21134
rect 470794 -1306 471414 20898
rect 470794 -1542 470826 -1306
rect 471062 -1542 471146 -1306
rect 471382 -1542 471414 -1306
rect 470794 -1626 471414 -1542
rect 470794 -1862 470826 -1626
rect 471062 -1862 471146 -1626
rect 471382 -1862 471414 -1626
rect 470794 -1894 471414 -1862
rect 471954 698614 472574 710042
rect 481954 711558 482574 711590
rect 481954 711322 481986 711558
rect 482222 711322 482306 711558
rect 482542 711322 482574 711558
rect 481954 711238 482574 711322
rect 481954 711002 481986 711238
rect 482222 711002 482306 711238
rect 482542 711002 482574 711238
rect 478234 709638 478854 709670
rect 478234 709402 478266 709638
rect 478502 709402 478586 709638
rect 478822 709402 478854 709638
rect 478234 709318 478854 709402
rect 478234 709082 478266 709318
rect 478502 709082 478586 709318
rect 478822 709082 478854 709318
rect 471954 698378 471986 698614
rect 472222 698378 472306 698614
rect 472542 698378 472574 698614
rect 471954 698294 472574 698378
rect 471954 698058 471986 698294
rect 472222 698058 472306 698294
rect 472542 698058 472574 698294
rect 471954 662614 472574 698058
rect 471954 662378 471986 662614
rect 472222 662378 472306 662614
rect 472542 662378 472574 662614
rect 471954 662294 472574 662378
rect 471954 662058 471986 662294
rect 472222 662058 472306 662294
rect 472542 662058 472574 662294
rect 471954 626614 472574 662058
rect 471954 626378 471986 626614
rect 472222 626378 472306 626614
rect 472542 626378 472574 626614
rect 471954 626294 472574 626378
rect 471954 626058 471986 626294
rect 472222 626058 472306 626294
rect 472542 626058 472574 626294
rect 471954 590614 472574 626058
rect 471954 590378 471986 590614
rect 472222 590378 472306 590614
rect 472542 590378 472574 590614
rect 471954 590294 472574 590378
rect 471954 590058 471986 590294
rect 472222 590058 472306 590294
rect 472542 590058 472574 590294
rect 471954 554614 472574 590058
rect 471954 554378 471986 554614
rect 472222 554378 472306 554614
rect 472542 554378 472574 554614
rect 471954 554294 472574 554378
rect 471954 554058 471986 554294
rect 472222 554058 472306 554294
rect 472542 554058 472574 554294
rect 471954 518614 472574 554058
rect 471954 518378 471986 518614
rect 472222 518378 472306 518614
rect 472542 518378 472574 518614
rect 471954 518294 472574 518378
rect 471954 518058 471986 518294
rect 472222 518058 472306 518294
rect 472542 518058 472574 518294
rect 471954 482614 472574 518058
rect 471954 482378 471986 482614
rect 472222 482378 472306 482614
rect 472542 482378 472574 482614
rect 471954 482294 472574 482378
rect 471954 482058 471986 482294
rect 472222 482058 472306 482294
rect 472542 482058 472574 482294
rect 471954 446614 472574 482058
rect 471954 446378 471986 446614
rect 472222 446378 472306 446614
rect 472542 446378 472574 446614
rect 471954 446294 472574 446378
rect 471954 446058 471986 446294
rect 472222 446058 472306 446294
rect 472542 446058 472574 446294
rect 471954 410614 472574 446058
rect 471954 410378 471986 410614
rect 472222 410378 472306 410614
rect 472542 410378 472574 410614
rect 471954 410294 472574 410378
rect 471954 410058 471986 410294
rect 472222 410058 472306 410294
rect 472542 410058 472574 410294
rect 471954 374614 472574 410058
rect 471954 374378 471986 374614
rect 472222 374378 472306 374614
rect 472542 374378 472574 374614
rect 471954 374294 472574 374378
rect 471954 374058 471986 374294
rect 472222 374058 472306 374294
rect 472542 374058 472574 374294
rect 471954 338614 472574 374058
rect 471954 338378 471986 338614
rect 472222 338378 472306 338614
rect 472542 338378 472574 338614
rect 471954 338294 472574 338378
rect 471954 338058 471986 338294
rect 472222 338058 472306 338294
rect 472542 338058 472574 338294
rect 471954 302614 472574 338058
rect 471954 302378 471986 302614
rect 472222 302378 472306 302614
rect 472542 302378 472574 302614
rect 471954 302294 472574 302378
rect 471954 302058 471986 302294
rect 472222 302058 472306 302294
rect 472542 302058 472574 302294
rect 471954 266614 472574 302058
rect 471954 266378 471986 266614
rect 472222 266378 472306 266614
rect 472542 266378 472574 266614
rect 471954 266294 472574 266378
rect 471954 266058 471986 266294
rect 472222 266058 472306 266294
rect 472542 266058 472574 266294
rect 471954 230614 472574 266058
rect 471954 230378 471986 230614
rect 472222 230378 472306 230614
rect 472542 230378 472574 230614
rect 471954 230294 472574 230378
rect 471954 230058 471986 230294
rect 472222 230058 472306 230294
rect 472542 230058 472574 230294
rect 471954 194614 472574 230058
rect 471954 194378 471986 194614
rect 472222 194378 472306 194614
rect 472542 194378 472574 194614
rect 471954 194294 472574 194378
rect 471954 194058 471986 194294
rect 472222 194058 472306 194294
rect 472542 194058 472574 194294
rect 471954 158614 472574 194058
rect 471954 158378 471986 158614
rect 472222 158378 472306 158614
rect 472542 158378 472574 158614
rect 471954 158294 472574 158378
rect 471954 158058 471986 158294
rect 472222 158058 472306 158294
rect 472542 158058 472574 158294
rect 471954 122614 472574 158058
rect 471954 122378 471986 122614
rect 472222 122378 472306 122614
rect 472542 122378 472574 122614
rect 471954 122294 472574 122378
rect 471954 122058 471986 122294
rect 472222 122058 472306 122294
rect 472542 122058 472574 122294
rect 471954 86614 472574 122058
rect 471954 86378 471986 86614
rect 472222 86378 472306 86614
rect 472542 86378 472574 86614
rect 471954 86294 472574 86378
rect 471954 86058 471986 86294
rect 472222 86058 472306 86294
rect 472542 86058 472574 86294
rect 471954 50614 472574 86058
rect 471954 50378 471986 50614
rect 472222 50378 472306 50614
rect 472542 50378 472574 50614
rect 471954 50294 472574 50378
rect 471954 50058 471986 50294
rect 472222 50058 472306 50294
rect 472542 50058 472574 50294
rect 471954 14614 472574 50058
rect 471954 14378 471986 14614
rect 472222 14378 472306 14614
rect 472542 14378 472574 14614
rect 471954 14294 472574 14378
rect 471954 14058 471986 14294
rect 472222 14058 472306 14294
rect 472542 14058 472574 14294
rect 468234 -4422 468266 -4186
rect 468502 -4422 468586 -4186
rect 468822 -4422 468854 -4186
rect 468234 -4506 468854 -4422
rect 468234 -4742 468266 -4506
rect 468502 -4742 468586 -4506
rect 468822 -4742 468854 -4506
rect 468234 -5734 468854 -4742
rect 461954 -7302 461986 -7066
rect 462222 -7302 462306 -7066
rect 462542 -7302 462574 -7066
rect 461954 -7386 462574 -7302
rect 461954 -7622 461986 -7386
rect 462222 -7622 462306 -7386
rect 462542 -7622 462574 -7386
rect 461954 -7654 462574 -7622
rect 471954 -6106 472574 14058
rect 474514 707718 475134 707750
rect 474514 707482 474546 707718
rect 474782 707482 474866 707718
rect 475102 707482 475134 707718
rect 474514 707398 475134 707482
rect 474514 707162 474546 707398
rect 474782 707162 474866 707398
rect 475102 707162 475134 707398
rect 474514 673174 475134 707162
rect 474514 672938 474546 673174
rect 474782 672938 474866 673174
rect 475102 672938 475134 673174
rect 474514 672854 475134 672938
rect 474514 672618 474546 672854
rect 474782 672618 474866 672854
rect 475102 672618 475134 672854
rect 474514 637174 475134 672618
rect 474514 636938 474546 637174
rect 474782 636938 474866 637174
rect 475102 636938 475134 637174
rect 474514 636854 475134 636938
rect 474514 636618 474546 636854
rect 474782 636618 474866 636854
rect 475102 636618 475134 636854
rect 474514 601174 475134 636618
rect 474514 600938 474546 601174
rect 474782 600938 474866 601174
rect 475102 600938 475134 601174
rect 474514 600854 475134 600938
rect 474514 600618 474546 600854
rect 474782 600618 474866 600854
rect 475102 600618 475134 600854
rect 474514 565174 475134 600618
rect 474514 564938 474546 565174
rect 474782 564938 474866 565174
rect 475102 564938 475134 565174
rect 474514 564854 475134 564938
rect 474514 564618 474546 564854
rect 474782 564618 474866 564854
rect 475102 564618 475134 564854
rect 474514 529174 475134 564618
rect 474514 528938 474546 529174
rect 474782 528938 474866 529174
rect 475102 528938 475134 529174
rect 474514 528854 475134 528938
rect 474514 528618 474546 528854
rect 474782 528618 474866 528854
rect 475102 528618 475134 528854
rect 474514 493174 475134 528618
rect 474514 492938 474546 493174
rect 474782 492938 474866 493174
rect 475102 492938 475134 493174
rect 474514 492854 475134 492938
rect 474514 492618 474546 492854
rect 474782 492618 474866 492854
rect 475102 492618 475134 492854
rect 474514 457174 475134 492618
rect 474514 456938 474546 457174
rect 474782 456938 474866 457174
rect 475102 456938 475134 457174
rect 474514 456854 475134 456938
rect 474514 456618 474546 456854
rect 474782 456618 474866 456854
rect 475102 456618 475134 456854
rect 474514 421174 475134 456618
rect 474514 420938 474546 421174
rect 474782 420938 474866 421174
rect 475102 420938 475134 421174
rect 474514 420854 475134 420938
rect 474514 420618 474546 420854
rect 474782 420618 474866 420854
rect 475102 420618 475134 420854
rect 474514 385174 475134 420618
rect 474514 384938 474546 385174
rect 474782 384938 474866 385174
rect 475102 384938 475134 385174
rect 474514 384854 475134 384938
rect 474514 384618 474546 384854
rect 474782 384618 474866 384854
rect 475102 384618 475134 384854
rect 474514 349174 475134 384618
rect 474514 348938 474546 349174
rect 474782 348938 474866 349174
rect 475102 348938 475134 349174
rect 474514 348854 475134 348938
rect 474514 348618 474546 348854
rect 474782 348618 474866 348854
rect 475102 348618 475134 348854
rect 474514 313174 475134 348618
rect 474514 312938 474546 313174
rect 474782 312938 474866 313174
rect 475102 312938 475134 313174
rect 474514 312854 475134 312938
rect 474514 312618 474546 312854
rect 474782 312618 474866 312854
rect 475102 312618 475134 312854
rect 474514 277174 475134 312618
rect 474514 276938 474546 277174
rect 474782 276938 474866 277174
rect 475102 276938 475134 277174
rect 474514 276854 475134 276938
rect 474514 276618 474546 276854
rect 474782 276618 474866 276854
rect 475102 276618 475134 276854
rect 474514 241174 475134 276618
rect 474514 240938 474546 241174
rect 474782 240938 474866 241174
rect 475102 240938 475134 241174
rect 474514 240854 475134 240938
rect 474514 240618 474546 240854
rect 474782 240618 474866 240854
rect 475102 240618 475134 240854
rect 474514 205174 475134 240618
rect 474514 204938 474546 205174
rect 474782 204938 474866 205174
rect 475102 204938 475134 205174
rect 474514 204854 475134 204938
rect 474514 204618 474546 204854
rect 474782 204618 474866 204854
rect 475102 204618 475134 204854
rect 474514 169174 475134 204618
rect 474514 168938 474546 169174
rect 474782 168938 474866 169174
rect 475102 168938 475134 169174
rect 474514 168854 475134 168938
rect 474514 168618 474546 168854
rect 474782 168618 474866 168854
rect 475102 168618 475134 168854
rect 474514 133174 475134 168618
rect 474514 132938 474546 133174
rect 474782 132938 474866 133174
rect 475102 132938 475134 133174
rect 474514 132854 475134 132938
rect 474514 132618 474546 132854
rect 474782 132618 474866 132854
rect 475102 132618 475134 132854
rect 474514 97174 475134 132618
rect 474514 96938 474546 97174
rect 474782 96938 474866 97174
rect 475102 96938 475134 97174
rect 474514 96854 475134 96938
rect 474514 96618 474546 96854
rect 474782 96618 474866 96854
rect 475102 96618 475134 96854
rect 474514 61174 475134 96618
rect 474514 60938 474546 61174
rect 474782 60938 474866 61174
rect 475102 60938 475134 61174
rect 474514 60854 475134 60938
rect 474514 60618 474546 60854
rect 474782 60618 474866 60854
rect 475102 60618 475134 60854
rect 474514 25174 475134 60618
rect 474514 24938 474546 25174
rect 474782 24938 474866 25174
rect 475102 24938 475134 25174
rect 474514 24854 475134 24938
rect 474514 24618 474546 24854
rect 474782 24618 474866 24854
rect 475102 24618 475134 24854
rect 474514 -3226 475134 24618
rect 474514 -3462 474546 -3226
rect 474782 -3462 474866 -3226
rect 475102 -3462 475134 -3226
rect 474514 -3546 475134 -3462
rect 474514 -3782 474546 -3546
rect 474782 -3782 474866 -3546
rect 475102 -3782 475134 -3546
rect 474514 -3814 475134 -3782
rect 478234 676894 478854 709082
rect 478234 676658 478266 676894
rect 478502 676658 478586 676894
rect 478822 676658 478854 676894
rect 478234 676574 478854 676658
rect 478234 676338 478266 676574
rect 478502 676338 478586 676574
rect 478822 676338 478854 676574
rect 478234 640894 478854 676338
rect 478234 640658 478266 640894
rect 478502 640658 478586 640894
rect 478822 640658 478854 640894
rect 478234 640574 478854 640658
rect 478234 640338 478266 640574
rect 478502 640338 478586 640574
rect 478822 640338 478854 640574
rect 478234 604894 478854 640338
rect 478234 604658 478266 604894
rect 478502 604658 478586 604894
rect 478822 604658 478854 604894
rect 478234 604574 478854 604658
rect 478234 604338 478266 604574
rect 478502 604338 478586 604574
rect 478822 604338 478854 604574
rect 478234 568894 478854 604338
rect 478234 568658 478266 568894
rect 478502 568658 478586 568894
rect 478822 568658 478854 568894
rect 478234 568574 478854 568658
rect 478234 568338 478266 568574
rect 478502 568338 478586 568574
rect 478822 568338 478854 568574
rect 478234 532894 478854 568338
rect 478234 532658 478266 532894
rect 478502 532658 478586 532894
rect 478822 532658 478854 532894
rect 478234 532574 478854 532658
rect 478234 532338 478266 532574
rect 478502 532338 478586 532574
rect 478822 532338 478854 532574
rect 478234 496894 478854 532338
rect 478234 496658 478266 496894
rect 478502 496658 478586 496894
rect 478822 496658 478854 496894
rect 478234 496574 478854 496658
rect 478234 496338 478266 496574
rect 478502 496338 478586 496574
rect 478822 496338 478854 496574
rect 478234 460894 478854 496338
rect 478234 460658 478266 460894
rect 478502 460658 478586 460894
rect 478822 460658 478854 460894
rect 478234 460574 478854 460658
rect 478234 460338 478266 460574
rect 478502 460338 478586 460574
rect 478822 460338 478854 460574
rect 478234 424894 478854 460338
rect 478234 424658 478266 424894
rect 478502 424658 478586 424894
rect 478822 424658 478854 424894
rect 478234 424574 478854 424658
rect 478234 424338 478266 424574
rect 478502 424338 478586 424574
rect 478822 424338 478854 424574
rect 478234 388894 478854 424338
rect 478234 388658 478266 388894
rect 478502 388658 478586 388894
rect 478822 388658 478854 388894
rect 478234 388574 478854 388658
rect 478234 388338 478266 388574
rect 478502 388338 478586 388574
rect 478822 388338 478854 388574
rect 478234 352894 478854 388338
rect 478234 352658 478266 352894
rect 478502 352658 478586 352894
rect 478822 352658 478854 352894
rect 478234 352574 478854 352658
rect 478234 352338 478266 352574
rect 478502 352338 478586 352574
rect 478822 352338 478854 352574
rect 478234 316894 478854 352338
rect 478234 316658 478266 316894
rect 478502 316658 478586 316894
rect 478822 316658 478854 316894
rect 478234 316574 478854 316658
rect 478234 316338 478266 316574
rect 478502 316338 478586 316574
rect 478822 316338 478854 316574
rect 478234 280894 478854 316338
rect 478234 280658 478266 280894
rect 478502 280658 478586 280894
rect 478822 280658 478854 280894
rect 478234 280574 478854 280658
rect 478234 280338 478266 280574
rect 478502 280338 478586 280574
rect 478822 280338 478854 280574
rect 478234 244894 478854 280338
rect 478234 244658 478266 244894
rect 478502 244658 478586 244894
rect 478822 244658 478854 244894
rect 478234 244574 478854 244658
rect 478234 244338 478266 244574
rect 478502 244338 478586 244574
rect 478822 244338 478854 244574
rect 478234 208894 478854 244338
rect 478234 208658 478266 208894
rect 478502 208658 478586 208894
rect 478822 208658 478854 208894
rect 478234 208574 478854 208658
rect 478234 208338 478266 208574
rect 478502 208338 478586 208574
rect 478822 208338 478854 208574
rect 478234 172894 478854 208338
rect 478234 172658 478266 172894
rect 478502 172658 478586 172894
rect 478822 172658 478854 172894
rect 478234 172574 478854 172658
rect 478234 172338 478266 172574
rect 478502 172338 478586 172574
rect 478822 172338 478854 172574
rect 478234 136894 478854 172338
rect 478234 136658 478266 136894
rect 478502 136658 478586 136894
rect 478822 136658 478854 136894
rect 478234 136574 478854 136658
rect 478234 136338 478266 136574
rect 478502 136338 478586 136574
rect 478822 136338 478854 136574
rect 478234 100894 478854 136338
rect 478234 100658 478266 100894
rect 478502 100658 478586 100894
rect 478822 100658 478854 100894
rect 478234 100574 478854 100658
rect 478234 100338 478266 100574
rect 478502 100338 478586 100574
rect 478822 100338 478854 100574
rect 478234 64894 478854 100338
rect 478234 64658 478266 64894
rect 478502 64658 478586 64894
rect 478822 64658 478854 64894
rect 478234 64574 478854 64658
rect 478234 64338 478266 64574
rect 478502 64338 478586 64574
rect 478822 64338 478854 64574
rect 478234 28894 478854 64338
rect 478234 28658 478266 28894
rect 478502 28658 478586 28894
rect 478822 28658 478854 28894
rect 478234 28574 478854 28658
rect 478234 28338 478266 28574
rect 478502 28338 478586 28574
rect 478822 28338 478854 28574
rect 478234 -5146 478854 28338
rect 480794 704838 481414 705830
rect 480794 704602 480826 704838
rect 481062 704602 481146 704838
rect 481382 704602 481414 704838
rect 480794 704518 481414 704602
rect 480794 704282 480826 704518
rect 481062 704282 481146 704518
rect 481382 704282 481414 704518
rect 480794 687454 481414 704282
rect 480794 687218 480826 687454
rect 481062 687218 481146 687454
rect 481382 687218 481414 687454
rect 480794 687134 481414 687218
rect 480794 686898 480826 687134
rect 481062 686898 481146 687134
rect 481382 686898 481414 687134
rect 480794 651454 481414 686898
rect 480794 651218 480826 651454
rect 481062 651218 481146 651454
rect 481382 651218 481414 651454
rect 480794 651134 481414 651218
rect 480794 650898 480826 651134
rect 481062 650898 481146 651134
rect 481382 650898 481414 651134
rect 480794 615454 481414 650898
rect 480794 615218 480826 615454
rect 481062 615218 481146 615454
rect 481382 615218 481414 615454
rect 480794 615134 481414 615218
rect 480794 614898 480826 615134
rect 481062 614898 481146 615134
rect 481382 614898 481414 615134
rect 480794 579454 481414 614898
rect 480794 579218 480826 579454
rect 481062 579218 481146 579454
rect 481382 579218 481414 579454
rect 480794 579134 481414 579218
rect 480794 578898 480826 579134
rect 481062 578898 481146 579134
rect 481382 578898 481414 579134
rect 480794 543454 481414 578898
rect 480794 543218 480826 543454
rect 481062 543218 481146 543454
rect 481382 543218 481414 543454
rect 480794 543134 481414 543218
rect 480794 542898 480826 543134
rect 481062 542898 481146 543134
rect 481382 542898 481414 543134
rect 480794 507454 481414 542898
rect 480794 507218 480826 507454
rect 481062 507218 481146 507454
rect 481382 507218 481414 507454
rect 480794 507134 481414 507218
rect 480794 506898 480826 507134
rect 481062 506898 481146 507134
rect 481382 506898 481414 507134
rect 480794 471454 481414 506898
rect 480794 471218 480826 471454
rect 481062 471218 481146 471454
rect 481382 471218 481414 471454
rect 480794 471134 481414 471218
rect 480794 470898 480826 471134
rect 481062 470898 481146 471134
rect 481382 470898 481414 471134
rect 480794 435454 481414 470898
rect 480794 435218 480826 435454
rect 481062 435218 481146 435454
rect 481382 435218 481414 435454
rect 480794 435134 481414 435218
rect 480794 434898 480826 435134
rect 481062 434898 481146 435134
rect 481382 434898 481414 435134
rect 480794 399454 481414 434898
rect 480794 399218 480826 399454
rect 481062 399218 481146 399454
rect 481382 399218 481414 399454
rect 480794 399134 481414 399218
rect 480794 398898 480826 399134
rect 481062 398898 481146 399134
rect 481382 398898 481414 399134
rect 480794 363454 481414 398898
rect 480794 363218 480826 363454
rect 481062 363218 481146 363454
rect 481382 363218 481414 363454
rect 480794 363134 481414 363218
rect 480794 362898 480826 363134
rect 481062 362898 481146 363134
rect 481382 362898 481414 363134
rect 480794 327454 481414 362898
rect 480794 327218 480826 327454
rect 481062 327218 481146 327454
rect 481382 327218 481414 327454
rect 480794 327134 481414 327218
rect 480794 326898 480826 327134
rect 481062 326898 481146 327134
rect 481382 326898 481414 327134
rect 480794 291454 481414 326898
rect 480794 291218 480826 291454
rect 481062 291218 481146 291454
rect 481382 291218 481414 291454
rect 480794 291134 481414 291218
rect 480794 290898 480826 291134
rect 481062 290898 481146 291134
rect 481382 290898 481414 291134
rect 480794 255454 481414 290898
rect 480794 255218 480826 255454
rect 481062 255218 481146 255454
rect 481382 255218 481414 255454
rect 480794 255134 481414 255218
rect 480794 254898 480826 255134
rect 481062 254898 481146 255134
rect 481382 254898 481414 255134
rect 480794 219454 481414 254898
rect 480794 219218 480826 219454
rect 481062 219218 481146 219454
rect 481382 219218 481414 219454
rect 480794 219134 481414 219218
rect 480794 218898 480826 219134
rect 481062 218898 481146 219134
rect 481382 218898 481414 219134
rect 480794 183454 481414 218898
rect 480794 183218 480826 183454
rect 481062 183218 481146 183454
rect 481382 183218 481414 183454
rect 480794 183134 481414 183218
rect 480794 182898 480826 183134
rect 481062 182898 481146 183134
rect 481382 182898 481414 183134
rect 480794 147454 481414 182898
rect 480794 147218 480826 147454
rect 481062 147218 481146 147454
rect 481382 147218 481414 147454
rect 480794 147134 481414 147218
rect 480794 146898 480826 147134
rect 481062 146898 481146 147134
rect 481382 146898 481414 147134
rect 480794 111454 481414 146898
rect 480794 111218 480826 111454
rect 481062 111218 481146 111454
rect 481382 111218 481414 111454
rect 480794 111134 481414 111218
rect 480794 110898 480826 111134
rect 481062 110898 481146 111134
rect 481382 110898 481414 111134
rect 480794 75454 481414 110898
rect 480794 75218 480826 75454
rect 481062 75218 481146 75454
rect 481382 75218 481414 75454
rect 480794 75134 481414 75218
rect 480794 74898 480826 75134
rect 481062 74898 481146 75134
rect 481382 74898 481414 75134
rect 480794 39454 481414 74898
rect 480794 39218 480826 39454
rect 481062 39218 481146 39454
rect 481382 39218 481414 39454
rect 480794 39134 481414 39218
rect 480794 38898 480826 39134
rect 481062 38898 481146 39134
rect 481382 38898 481414 39134
rect 480794 3454 481414 38898
rect 480794 3218 480826 3454
rect 481062 3218 481146 3454
rect 481382 3218 481414 3454
rect 480794 3134 481414 3218
rect 480794 2898 480826 3134
rect 481062 2898 481146 3134
rect 481382 2898 481414 3134
rect 480794 -346 481414 2898
rect 480794 -582 480826 -346
rect 481062 -582 481146 -346
rect 481382 -582 481414 -346
rect 480794 -666 481414 -582
rect 480794 -902 480826 -666
rect 481062 -902 481146 -666
rect 481382 -902 481414 -666
rect 480794 -1894 481414 -902
rect 481954 680614 482574 711002
rect 491954 710598 492574 711590
rect 491954 710362 491986 710598
rect 492222 710362 492306 710598
rect 492542 710362 492574 710598
rect 491954 710278 492574 710362
rect 491954 710042 491986 710278
rect 492222 710042 492306 710278
rect 492542 710042 492574 710278
rect 488234 708678 488854 709670
rect 488234 708442 488266 708678
rect 488502 708442 488586 708678
rect 488822 708442 488854 708678
rect 488234 708358 488854 708442
rect 488234 708122 488266 708358
rect 488502 708122 488586 708358
rect 488822 708122 488854 708358
rect 481954 680378 481986 680614
rect 482222 680378 482306 680614
rect 482542 680378 482574 680614
rect 481954 680294 482574 680378
rect 481954 680058 481986 680294
rect 482222 680058 482306 680294
rect 482542 680058 482574 680294
rect 481954 644614 482574 680058
rect 481954 644378 481986 644614
rect 482222 644378 482306 644614
rect 482542 644378 482574 644614
rect 481954 644294 482574 644378
rect 481954 644058 481986 644294
rect 482222 644058 482306 644294
rect 482542 644058 482574 644294
rect 481954 608614 482574 644058
rect 481954 608378 481986 608614
rect 482222 608378 482306 608614
rect 482542 608378 482574 608614
rect 481954 608294 482574 608378
rect 481954 608058 481986 608294
rect 482222 608058 482306 608294
rect 482542 608058 482574 608294
rect 481954 572614 482574 608058
rect 481954 572378 481986 572614
rect 482222 572378 482306 572614
rect 482542 572378 482574 572614
rect 481954 572294 482574 572378
rect 481954 572058 481986 572294
rect 482222 572058 482306 572294
rect 482542 572058 482574 572294
rect 481954 536614 482574 572058
rect 481954 536378 481986 536614
rect 482222 536378 482306 536614
rect 482542 536378 482574 536614
rect 481954 536294 482574 536378
rect 481954 536058 481986 536294
rect 482222 536058 482306 536294
rect 482542 536058 482574 536294
rect 481954 500614 482574 536058
rect 481954 500378 481986 500614
rect 482222 500378 482306 500614
rect 482542 500378 482574 500614
rect 481954 500294 482574 500378
rect 481954 500058 481986 500294
rect 482222 500058 482306 500294
rect 482542 500058 482574 500294
rect 481954 464614 482574 500058
rect 481954 464378 481986 464614
rect 482222 464378 482306 464614
rect 482542 464378 482574 464614
rect 481954 464294 482574 464378
rect 481954 464058 481986 464294
rect 482222 464058 482306 464294
rect 482542 464058 482574 464294
rect 481954 428614 482574 464058
rect 481954 428378 481986 428614
rect 482222 428378 482306 428614
rect 482542 428378 482574 428614
rect 481954 428294 482574 428378
rect 481954 428058 481986 428294
rect 482222 428058 482306 428294
rect 482542 428058 482574 428294
rect 481954 392614 482574 428058
rect 481954 392378 481986 392614
rect 482222 392378 482306 392614
rect 482542 392378 482574 392614
rect 481954 392294 482574 392378
rect 481954 392058 481986 392294
rect 482222 392058 482306 392294
rect 482542 392058 482574 392294
rect 481954 356614 482574 392058
rect 481954 356378 481986 356614
rect 482222 356378 482306 356614
rect 482542 356378 482574 356614
rect 481954 356294 482574 356378
rect 481954 356058 481986 356294
rect 482222 356058 482306 356294
rect 482542 356058 482574 356294
rect 481954 320614 482574 356058
rect 481954 320378 481986 320614
rect 482222 320378 482306 320614
rect 482542 320378 482574 320614
rect 481954 320294 482574 320378
rect 481954 320058 481986 320294
rect 482222 320058 482306 320294
rect 482542 320058 482574 320294
rect 481954 284614 482574 320058
rect 481954 284378 481986 284614
rect 482222 284378 482306 284614
rect 482542 284378 482574 284614
rect 481954 284294 482574 284378
rect 481954 284058 481986 284294
rect 482222 284058 482306 284294
rect 482542 284058 482574 284294
rect 481954 248614 482574 284058
rect 481954 248378 481986 248614
rect 482222 248378 482306 248614
rect 482542 248378 482574 248614
rect 481954 248294 482574 248378
rect 481954 248058 481986 248294
rect 482222 248058 482306 248294
rect 482542 248058 482574 248294
rect 481954 212614 482574 248058
rect 481954 212378 481986 212614
rect 482222 212378 482306 212614
rect 482542 212378 482574 212614
rect 481954 212294 482574 212378
rect 481954 212058 481986 212294
rect 482222 212058 482306 212294
rect 482542 212058 482574 212294
rect 481954 176614 482574 212058
rect 481954 176378 481986 176614
rect 482222 176378 482306 176614
rect 482542 176378 482574 176614
rect 481954 176294 482574 176378
rect 481954 176058 481986 176294
rect 482222 176058 482306 176294
rect 482542 176058 482574 176294
rect 481954 140614 482574 176058
rect 481954 140378 481986 140614
rect 482222 140378 482306 140614
rect 482542 140378 482574 140614
rect 481954 140294 482574 140378
rect 481954 140058 481986 140294
rect 482222 140058 482306 140294
rect 482542 140058 482574 140294
rect 481954 104614 482574 140058
rect 481954 104378 481986 104614
rect 482222 104378 482306 104614
rect 482542 104378 482574 104614
rect 481954 104294 482574 104378
rect 481954 104058 481986 104294
rect 482222 104058 482306 104294
rect 482542 104058 482574 104294
rect 481954 68614 482574 104058
rect 481954 68378 481986 68614
rect 482222 68378 482306 68614
rect 482542 68378 482574 68614
rect 481954 68294 482574 68378
rect 481954 68058 481986 68294
rect 482222 68058 482306 68294
rect 482542 68058 482574 68294
rect 481954 32614 482574 68058
rect 481954 32378 481986 32614
rect 482222 32378 482306 32614
rect 482542 32378 482574 32614
rect 481954 32294 482574 32378
rect 481954 32058 481986 32294
rect 482222 32058 482306 32294
rect 482542 32058 482574 32294
rect 478234 -5382 478266 -5146
rect 478502 -5382 478586 -5146
rect 478822 -5382 478854 -5146
rect 478234 -5466 478854 -5382
rect 478234 -5702 478266 -5466
rect 478502 -5702 478586 -5466
rect 478822 -5702 478854 -5466
rect 478234 -5734 478854 -5702
rect 471954 -6342 471986 -6106
rect 472222 -6342 472306 -6106
rect 472542 -6342 472574 -6106
rect 471954 -6426 472574 -6342
rect 471954 -6662 471986 -6426
rect 472222 -6662 472306 -6426
rect 472542 -6662 472574 -6426
rect 471954 -7654 472574 -6662
rect 481954 -7066 482574 32058
rect 484514 706758 485134 707750
rect 484514 706522 484546 706758
rect 484782 706522 484866 706758
rect 485102 706522 485134 706758
rect 484514 706438 485134 706522
rect 484514 706202 484546 706438
rect 484782 706202 484866 706438
rect 485102 706202 485134 706438
rect 484514 691174 485134 706202
rect 484514 690938 484546 691174
rect 484782 690938 484866 691174
rect 485102 690938 485134 691174
rect 484514 690854 485134 690938
rect 484514 690618 484546 690854
rect 484782 690618 484866 690854
rect 485102 690618 485134 690854
rect 484514 655174 485134 690618
rect 484514 654938 484546 655174
rect 484782 654938 484866 655174
rect 485102 654938 485134 655174
rect 484514 654854 485134 654938
rect 484514 654618 484546 654854
rect 484782 654618 484866 654854
rect 485102 654618 485134 654854
rect 484514 619174 485134 654618
rect 484514 618938 484546 619174
rect 484782 618938 484866 619174
rect 485102 618938 485134 619174
rect 484514 618854 485134 618938
rect 484514 618618 484546 618854
rect 484782 618618 484866 618854
rect 485102 618618 485134 618854
rect 484514 583174 485134 618618
rect 484514 582938 484546 583174
rect 484782 582938 484866 583174
rect 485102 582938 485134 583174
rect 484514 582854 485134 582938
rect 484514 582618 484546 582854
rect 484782 582618 484866 582854
rect 485102 582618 485134 582854
rect 484514 547174 485134 582618
rect 484514 546938 484546 547174
rect 484782 546938 484866 547174
rect 485102 546938 485134 547174
rect 484514 546854 485134 546938
rect 484514 546618 484546 546854
rect 484782 546618 484866 546854
rect 485102 546618 485134 546854
rect 484514 511174 485134 546618
rect 484514 510938 484546 511174
rect 484782 510938 484866 511174
rect 485102 510938 485134 511174
rect 484514 510854 485134 510938
rect 484514 510618 484546 510854
rect 484782 510618 484866 510854
rect 485102 510618 485134 510854
rect 484514 475174 485134 510618
rect 484514 474938 484546 475174
rect 484782 474938 484866 475174
rect 485102 474938 485134 475174
rect 484514 474854 485134 474938
rect 484514 474618 484546 474854
rect 484782 474618 484866 474854
rect 485102 474618 485134 474854
rect 484514 439174 485134 474618
rect 484514 438938 484546 439174
rect 484782 438938 484866 439174
rect 485102 438938 485134 439174
rect 484514 438854 485134 438938
rect 484514 438618 484546 438854
rect 484782 438618 484866 438854
rect 485102 438618 485134 438854
rect 484514 403174 485134 438618
rect 484514 402938 484546 403174
rect 484782 402938 484866 403174
rect 485102 402938 485134 403174
rect 484514 402854 485134 402938
rect 484514 402618 484546 402854
rect 484782 402618 484866 402854
rect 485102 402618 485134 402854
rect 484514 367174 485134 402618
rect 484514 366938 484546 367174
rect 484782 366938 484866 367174
rect 485102 366938 485134 367174
rect 484514 366854 485134 366938
rect 484514 366618 484546 366854
rect 484782 366618 484866 366854
rect 485102 366618 485134 366854
rect 484514 331174 485134 366618
rect 484514 330938 484546 331174
rect 484782 330938 484866 331174
rect 485102 330938 485134 331174
rect 484514 330854 485134 330938
rect 484514 330618 484546 330854
rect 484782 330618 484866 330854
rect 485102 330618 485134 330854
rect 484514 295174 485134 330618
rect 484514 294938 484546 295174
rect 484782 294938 484866 295174
rect 485102 294938 485134 295174
rect 484514 294854 485134 294938
rect 484514 294618 484546 294854
rect 484782 294618 484866 294854
rect 485102 294618 485134 294854
rect 484514 259174 485134 294618
rect 484514 258938 484546 259174
rect 484782 258938 484866 259174
rect 485102 258938 485134 259174
rect 484514 258854 485134 258938
rect 484514 258618 484546 258854
rect 484782 258618 484866 258854
rect 485102 258618 485134 258854
rect 484514 223174 485134 258618
rect 484514 222938 484546 223174
rect 484782 222938 484866 223174
rect 485102 222938 485134 223174
rect 484514 222854 485134 222938
rect 484514 222618 484546 222854
rect 484782 222618 484866 222854
rect 485102 222618 485134 222854
rect 484514 187174 485134 222618
rect 484514 186938 484546 187174
rect 484782 186938 484866 187174
rect 485102 186938 485134 187174
rect 484514 186854 485134 186938
rect 484514 186618 484546 186854
rect 484782 186618 484866 186854
rect 485102 186618 485134 186854
rect 484514 151174 485134 186618
rect 484514 150938 484546 151174
rect 484782 150938 484866 151174
rect 485102 150938 485134 151174
rect 484514 150854 485134 150938
rect 484514 150618 484546 150854
rect 484782 150618 484866 150854
rect 485102 150618 485134 150854
rect 484514 115174 485134 150618
rect 484514 114938 484546 115174
rect 484782 114938 484866 115174
rect 485102 114938 485134 115174
rect 484514 114854 485134 114938
rect 484514 114618 484546 114854
rect 484782 114618 484866 114854
rect 485102 114618 485134 114854
rect 484514 79174 485134 114618
rect 484514 78938 484546 79174
rect 484782 78938 484866 79174
rect 485102 78938 485134 79174
rect 484514 78854 485134 78938
rect 484514 78618 484546 78854
rect 484782 78618 484866 78854
rect 485102 78618 485134 78854
rect 484514 43174 485134 78618
rect 484514 42938 484546 43174
rect 484782 42938 484866 43174
rect 485102 42938 485134 43174
rect 484514 42854 485134 42938
rect 484514 42618 484546 42854
rect 484782 42618 484866 42854
rect 485102 42618 485134 42854
rect 484514 7174 485134 42618
rect 484514 6938 484546 7174
rect 484782 6938 484866 7174
rect 485102 6938 485134 7174
rect 484514 6854 485134 6938
rect 484514 6618 484546 6854
rect 484782 6618 484866 6854
rect 485102 6618 485134 6854
rect 484514 -2266 485134 6618
rect 484514 -2502 484546 -2266
rect 484782 -2502 484866 -2266
rect 485102 -2502 485134 -2266
rect 484514 -2586 485134 -2502
rect 484514 -2822 484546 -2586
rect 484782 -2822 484866 -2586
rect 485102 -2822 485134 -2586
rect 484514 -3814 485134 -2822
rect 488234 694894 488854 708122
rect 488234 694658 488266 694894
rect 488502 694658 488586 694894
rect 488822 694658 488854 694894
rect 488234 694574 488854 694658
rect 488234 694338 488266 694574
rect 488502 694338 488586 694574
rect 488822 694338 488854 694574
rect 488234 658894 488854 694338
rect 488234 658658 488266 658894
rect 488502 658658 488586 658894
rect 488822 658658 488854 658894
rect 488234 658574 488854 658658
rect 488234 658338 488266 658574
rect 488502 658338 488586 658574
rect 488822 658338 488854 658574
rect 488234 622894 488854 658338
rect 488234 622658 488266 622894
rect 488502 622658 488586 622894
rect 488822 622658 488854 622894
rect 488234 622574 488854 622658
rect 488234 622338 488266 622574
rect 488502 622338 488586 622574
rect 488822 622338 488854 622574
rect 488234 586894 488854 622338
rect 488234 586658 488266 586894
rect 488502 586658 488586 586894
rect 488822 586658 488854 586894
rect 488234 586574 488854 586658
rect 488234 586338 488266 586574
rect 488502 586338 488586 586574
rect 488822 586338 488854 586574
rect 488234 550894 488854 586338
rect 488234 550658 488266 550894
rect 488502 550658 488586 550894
rect 488822 550658 488854 550894
rect 488234 550574 488854 550658
rect 488234 550338 488266 550574
rect 488502 550338 488586 550574
rect 488822 550338 488854 550574
rect 488234 514894 488854 550338
rect 488234 514658 488266 514894
rect 488502 514658 488586 514894
rect 488822 514658 488854 514894
rect 488234 514574 488854 514658
rect 488234 514338 488266 514574
rect 488502 514338 488586 514574
rect 488822 514338 488854 514574
rect 488234 478894 488854 514338
rect 488234 478658 488266 478894
rect 488502 478658 488586 478894
rect 488822 478658 488854 478894
rect 488234 478574 488854 478658
rect 488234 478338 488266 478574
rect 488502 478338 488586 478574
rect 488822 478338 488854 478574
rect 488234 442894 488854 478338
rect 488234 442658 488266 442894
rect 488502 442658 488586 442894
rect 488822 442658 488854 442894
rect 488234 442574 488854 442658
rect 488234 442338 488266 442574
rect 488502 442338 488586 442574
rect 488822 442338 488854 442574
rect 488234 406894 488854 442338
rect 488234 406658 488266 406894
rect 488502 406658 488586 406894
rect 488822 406658 488854 406894
rect 488234 406574 488854 406658
rect 488234 406338 488266 406574
rect 488502 406338 488586 406574
rect 488822 406338 488854 406574
rect 488234 370894 488854 406338
rect 488234 370658 488266 370894
rect 488502 370658 488586 370894
rect 488822 370658 488854 370894
rect 488234 370574 488854 370658
rect 488234 370338 488266 370574
rect 488502 370338 488586 370574
rect 488822 370338 488854 370574
rect 488234 334894 488854 370338
rect 488234 334658 488266 334894
rect 488502 334658 488586 334894
rect 488822 334658 488854 334894
rect 488234 334574 488854 334658
rect 488234 334338 488266 334574
rect 488502 334338 488586 334574
rect 488822 334338 488854 334574
rect 488234 298894 488854 334338
rect 488234 298658 488266 298894
rect 488502 298658 488586 298894
rect 488822 298658 488854 298894
rect 488234 298574 488854 298658
rect 488234 298338 488266 298574
rect 488502 298338 488586 298574
rect 488822 298338 488854 298574
rect 488234 262894 488854 298338
rect 488234 262658 488266 262894
rect 488502 262658 488586 262894
rect 488822 262658 488854 262894
rect 488234 262574 488854 262658
rect 488234 262338 488266 262574
rect 488502 262338 488586 262574
rect 488822 262338 488854 262574
rect 488234 226894 488854 262338
rect 488234 226658 488266 226894
rect 488502 226658 488586 226894
rect 488822 226658 488854 226894
rect 488234 226574 488854 226658
rect 488234 226338 488266 226574
rect 488502 226338 488586 226574
rect 488822 226338 488854 226574
rect 488234 190894 488854 226338
rect 488234 190658 488266 190894
rect 488502 190658 488586 190894
rect 488822 190658 488854 190894
rect 488234 190574 488854 190658
rect 488234 190338 488266 190574
rect 488502 190338 488586 190574
rect 488822 190338 488854 190574
rect 488234 154894 488854 190338
rect 488234 154658 488266 154894
rect 488502 154658 488586 154894
rect 488822 154658 488854 154894
rect 488234 154574 488854 154658
rect 488234 154338 488266 154574
rect 488502 154338 488586 154574
rect 488822 154338 488854 154574
rect 488234 118894 488854 154338
rect 488234 118658 488266 118894
rect 488502 118658 488586 118894
rect 488822 118658 488854 118894
rect 488234 118574 488854 118658
rect 488234 118338 488266 118574
rect 488502 118338 488586 118574
rect 488822 118338 488854 118574
rect 488234 82894 488854 118338
rect 488234 82658 488266 82894
rect 488502 82658 488586 82894
rect 488822 82658 488854 82894
rect 488234 82574 488854 82658
rect 488234 82338 488266 82574
rect 488502 82338 488586 82574
rect 488822 82338 488854 82574
rect 488234 46894 488854 82338
rect 488234 46658 488266 46894
rect 488502 46658 488586 46894
rect 488822 46658 488854 46894
rect 488234 46574 488854 46658
rect 488234 46338 488266 46574
rect 488502 46338 488586 46574
rect 488822 46338 488854 46574
rect 488234 10894 488854 46338
rect 488234 10658 488266 10894
rect 488502 10658 488586 10894
rect 488822 10658 488854 10894
rect 488234 10574 488854 10658
rect 488234 10338 488266 10574
rect 488502 10338 488586 10574
rect 488822 10338 488854 10574
rect 488234 -4186 488854 10338
rect 490794 705798 491414 705830
rect 490794 705562 490826 705798
rect 491062 705562 491146 705798
rect 491382 705562 491414 705798
rect 490794 705478 491414 705562
rect 490794 705242 490826 705478
rect 491062 705242 491146 705478
rect 491382 705242 491414 705478
rect 490794 669454 491414 705242
rect 490794 669218 490826 669454
rect 491062 669218 491146 669454
rect 491382 669218 491414 669454
rect 490794 669134 491414 669218
rect 490794 668898 490826 669134
rect 491062 668898 491146 669134
rect 491382 668898 491414 669134
rect 490794 633454 491414 668898
rect 490794 633218 490826 633454
rect 491062 633218 491146 633454
rect 491382 633218 491414 633454
rect 490794 633134 491414 633218
rect 490794 632898 490826 633134
rect 491062 632898 491146 633134
rect 491382 632898 491414 633134
rect 490794 597454 491414 632898
rect 490794 597218 490826 597454
rect 491062 597218 491146 597454
rect 491382 597218 491414 597454
rect 490794 597134 491414 597218
rect 490794 596898 490826 597134
rect 491062 596898 491146 597134
rect 491382 596898 491414 597134
rect 490794 561454 491414 596898
rect 490794 561218 490826 561454
rect 491062 561218 491146 561454
rect 491382 561218 491414 561454
rect 490794 561134 491414 561218
rect 490794 560898 490826 561134
rect 491062 560898 491146 561134
rect 491382 560898 491414 561134
rect 490794 525454 491414 560898
rect 490794 525218 490826 525454
rect 491062 525218 491146 525454
rect 491382 525218 491414 525454
rect 490794 525134 491414 525218
rect 490794 524898 490826 525134
rect 491062 524898 491146 525134
rect 491382 524898 491414 525134
rect 490794 489454 491414 524898
rect 490794 489218 490826 489454
rect 491062 489218 491146 489454
rect 491382 489218 491414 489454
rect 490794 489134 491414 489218
rect 490794 488898 490826 489134
rect 491062 488898 491146 489134
rect 491382 488898 491414 489134
rect 490794 453454 491414 488898
rect 490794 453218 490826 453454
rect 491062 453218 491146 453454
rect 491382 453218 491414 453454
rect 490794 453134 491414 453218
rect 490794 452898 490826 453134
rect 491062 452898 491146 453134
rect 491382 452898 491414 453134
rect 490794 417454 491414 452898
rect 490794 417218 490826 417454
rect 491062 417218 491146 417454
rect 491382 417218 491414 417454
rect 490794 417134 491414 417218
rect 490794 416898 490826 417134
rect 491062 416898 491146 417134
rect 491382 416898 491414 417134
rect 490794 381454 491414 416898
rect 490794 381218 490826 381454
rect 491062 381218 491146 381454
rect 491382 381218 491414 381454
rect 490794 381134 491414 381218
rect 490794 380898 490826 381134
rect 491062 380898 491146 381134
rect 491382 380898 491414 381134
rect 490794 345454 491414 380898
rect 490794 345218 490826 345454
rect 491062 345218 491146 345454
rect 491382 345218 491414 345454
rect 490794 345134 491414 345218
rect 490794 344898 490826 345134
rect 491062 344898 491146 345134
rect 491382 344898 491414 345134
rect 490794 309454 491414 344898
rect 490794 309218 490826 309454
rect 491062 309218 491146 309454
rect 491382 309218 491414 309454
rect 490794 309134 491414 309218
rect 490794 308898 490826 309134
rect 491062 308898 491146 309134
rect 491382 308898 491414 309134
rect 490794 273454 491414 308898
rect 490794 273218 490826 273454
rect 491062 273218 491146 273454
rect 491382 273218 491414 273454
rect 490794 273134 491414 273218
rect 490794 272898 490826 273134
rect 491062 272898 491146 273134
rect 491382 272898 491414 273134
rect 490794 237454 491414 272898
rect 490794 237218 490826 237454
rect 491062 237218 491146 237454
rect 491382 237218 491414 237454
rect 490794 237134 491414 237218
rect 490794 236898 490826 237134
rect 491062 236898 491146 237134
rect 491382 236898 491414 237134
rect 490794 201454 491414 236898
rect 490794 201218 490826 201454
rect 491062 201218 491146 201454
rect 491382 201218 491414 201454
rect 490794 201134 491414 201218
rect 490794 200898 490826 201134
rect 491062 200898 491146 201134
rect 491382 200898 491414 201134
rect 490794 165454 491414 200898
rect 490794 165218 490826 165454
rect 491062 165218 491146 165454
rect 491382 165218 491414 165454
rect 490794 165134 491414 165218
rect 490794 164898 490826 165134
rect 491062 164898 491146 165134
rect 491382 164898 491414 165134
rect 490794 129454 491414 164898
rect 490794 129218 490826 129454
rect 491062 129218 491146 129454
rect 491382 129218 491414 129454
rect 490794 129134 491414 129218
rect 490794 128898 490826 129134
rect 491062 128898 491146 129134
rect 491382 128898 491414 129134
rect 490794 93454 491414 128898
rect 490794 93218 490826 93454
rect 491062 93218 491146 93454
rect 491382 93218 491414 93454
rect 490794 93134 491414 93218
rect 490794 92898 490826 93134
rect 491062 92898 491146 93134
rect 491382 92898 491414 93134
rect 490794 57454 491414 92898
rect 490794 57218 490826 57454
rect 491062 57218 491146 57454
rect 491382 57218 491414 57454
rect 490794 57134 491414 57218
rect 490794 56898 490826 57134
rect 491062 56898 491146 57134
rect 491382 56898 491414 57134
rect 490794 21454 491414 56898
rect 490794 21218 490826 21454
rect 491062 21218 491146 21454
rect 491382 21218 491414 21454
rect 490794 21134 491414 21218
rect 490794 20898 490826 21134
rect 491062 20898 491146 21134
rect 491382 20898 491414 21134
rect 490794 -1306 491414 20898
rect 490794 -1542 490826 -1306
rect 491062 -1542 491146 -1306
rect 491382 -1542 491414 -1306
rect 490794 -1626 491414 -1542
rect 490794 -1862 490826 -1626
rect 491062 -1862 491146 -1626
rect 491382 -1862 491414 -1626
rect 490794 -1894 491414 -1862
rect 491954 698614 492574 710042
rect 501954 711558 502574 711590
rect 501954 711322 501986 711558
rect 502222 711322 502306 711558
rect 502542 711322 502574 711558
rect 501954 711238 502574 711322
rect 501954 711002 501986 711238
rect 502222 711002 502306 711238
rect 502542 711002 502574 711238
rect 498234 709638 498854 709670
rect 498234 709402 498266 709638
rect 498502 709402 498586 709638
rect 498822 709402 498854 709638
rect 498234 709318 498854 709402
rect 498234 709082 498266 709318
rect 498502 709082 498586 709318
rect 498822 709082 498854 709318
rect 491954 698378 491986 698614
rect 492222 698378 492306 698614
rect 492542 698378 492574 698614
rect 491954 698294 492574 698378
rect 491954 698058 491986 698294
rect 492222 698058 492306 698294
rect 492542 698058 492574 698294
rect 491954 662614 492574 698058
rect 491954 662378 491986 662614
rect 492222 662378 492306 662614
rect 492542 662378 492574 662614
rect 491954 662294 492574 662378
rect 491954 662058 491986 662294
rect 492222 662058 492306 662294
rect 492542 662058 492574 662294
rect 491954 626614 492574 662058
rect 491954 626378 491986 626614
rect 492222 626378 492306 626614
rect 492542 626378 492574 626614
rect 491954 626294 492574 626378
rect 491954 626058 491986 626294
rect 492222 626058 492306 626294
rect 492542 626058 492574 626294
rect 491954 590614 492574 626058
rect 491954 590378 491986 590614
rect 492222 590378 492306 590614
rect 492542 590378 492574 590614
rect 491954 590294 492574 590378
rect 491954 590058 491986 590294
rect 492222 590058 492306 590294
rect 492542 590058 492574 590294
rect 491954 554614 492574 590058
rect 491954 554378 491986 554614
rect 492222 554378 492306 554614
rect 492542 554378 492574 554614
rect 491954 554294 492574 554378
rect 491954 554058 491986 554294
rect 492222 554058 492306 554294
rect 492542 554058 492574 554294
rect 491954 518614 492574 554058
rect 491954 518378 491986 518614
rect 492222 518378 492306 518614
rect 492542 518378 492574 518614
rect 491954 518294 492574 518378
rect 491954 518058 491986 518294
rect 492222 518058 492306 518294
rect 492542 518058 492574 518294
rect 491954 482614 492574 518058
rect 491954 482378 491986 482614
rect 492222 482378 492306 482614
rect 492542 482378 492574 482614
rect 491954 482294 492574 482378
rect 491954 482058 491986 482294
rect 492222 482058 492306 482294
rect 492542 482058 492574 482294
rect 491954 446614 492574 482058
rect 491954 446378 491986 446614
rect 492222 446378 492306 446614
rect 492542 446378 492574 446614
rect 491954 446294 492574 446378
rect 491954 446058 491986 446294
rect 492222 446058 492306 446294
rect 492542 446058 492574 446294
rect 491954 410614 492574 446058
rect 491954 410378 491986 410614
rect 492222 410378 492306 410614
rect 492542 410378 492574 410614
rect 491954 410294 492574 410378
rect 491954 410058 491986 410294
rect 492222 410058 492306 410294
rect 492542 410058 492574 410294
rect 491954 374614 492574 410058
rect 491954 374378 491986 374614
rect 492222 374378 492306 374614
rect 492542 374378 492574 374614
rect 491954 374294 492574 374378
rect 491954 374058 491986 374294
rect 492222 374058 492306 374294
rect 492542 374058 492574 374294
rect 491954 338614 492574 374058
rect 491954 338378 491986 338614
rect 492222 338378 492306 338614
rect 492542 338378 492574 338614
rect 491954 338294 492574 338378
rect 491954 338058 491986 338294
rect 492222 338058 492306 338294
rect 492542 338058 492574 338294
rect 491954 302614 492574 338058
rect 491954 302378 491986 302614
rect 492222 302378 492306 302614
rect 492542 302378 492574 302614
rect 491954 302294 492574 302378
rect 491954 302058 491986 302294
rect 492222 302058 492306 302294
rect 492542 302058 492574 302294
rect 491954 266614 492574 302058
rect 491954 266378 491986 266614
rect 492222 266378 492306 266614
rect 492542 266378 492574 266614
rect 491954 266294 492574 266378
rect 491954 266058 491986 266294
rect 492222 266058 492306 266294
rect 492542 266058 492574 266294
rect 491954 230614 492574 266058
rect 491954 230378 491986 230614
rect 492222 230378 492306 230614
rect 492542 230378 492574 230614
rect 491954 230294 492574 230378
rect 491954 230058 491986 230294
rect 492222 230058 492306 230294
rect 492542 230058 492574 230294
rect 491954 194614 492574 230058
rect 491954 194378 491986 194614
rect 492222 194378 492306 194614
rect 492542 194378 492574 194614
rect 491954 194294 492574 194378
rect 491954 194058 491986 194294
rect 492222 194058 492306 194294
rect 492542 194058 492574 194294
rect 491954 158614 492574 194058
rect 491954 158378 491986 158614
rect 492222 158378 492306 158614
rect 492542 158378 492574 158614
rect 491954 158294 492574 158378
rect 491954 158058 491986 158294
rect 492222 158058 492306 158294
rect 492542 158058 492574 158294
rect 491954 122614 492574 158058
rect 491954 122378 491986 122614
rect 492222 122378 492306 122614
rect 492542 122378 492574 122614
rect 491954 122294 492574 122378
rect 491954 122058 491986 122294
rect 492222 122058 492306 122294
rect 492542 122058 492574 122294
rect 491954 86614 492574 122058
rect 491954 86378 491986 86614
rect 492222 86378 492306 86614
rect 492542 86378 492574 86614
rect 491954 86294 492574 86378
rect 491954 86058 491986 86294
rect 492222 86058 492306 86294
rect 492542 86058 492574 86294
rect 491954 50614 492574 86058
rect 491954 50378 491986 50614
rect 492222 50378 492306 50614
rect 492542 50378 492574 50614
rect 491954 50294 492574 50378
rect 491954 50058 491986 50294
rect 492222 50058 492306 50294
rect 492542 50058 492574 50294
rect 491954 14614 492574 50058
rect 491954 14378 491986 14614
rect 492222 14378 492306 14614
rect 492542 14378 492574 14614
rect 491954 14294 492574 14378
rect 491954 14058 491986 14294
rect 492222 14058 492306 14294
rect 492542 14058 492574 14294
rect 488234 -4422 488266 -4186
rect 488502 -4422 488586 -4186
rect 488822 -4422 488854 -4186
rect 488234 -4506 488854 -4422
rect 488234 -4742 488266 -4506
rect 488502 -4742 488586 -4506
rect 488822 -4742 488854 -4506
rect 488234 -5734 488854 -4742
rect 481954 -7302 481986 -7066
rect 482222 -7302 482306 -7066
rect 482542 -7302 482574 -7066
rect 481954 -7386 482574 -7302
rect 481954 -7622 481986 -7386
rect 482222 -7622 482306 -7386
rect 482542 -7622 482574 -7386
rect 481954 -7654 482574 -7622
rect 491954 -6106 492574 14058
rect 494514 707718 495134 707750
rect 494514 707482 494546 707718
rect 494782 707482 494866 707718
rect 495102 707482 495134 707718
rect 494514 707398 495134 707482
rect 494514 707162 494546 707398
rect 494782 707162 494866 707398
rect 495102 707162 495134 707398
rect 494514 673174 495134 707162
rect 494514 672938 494546 673174
rect 494782 672938 494866 673174
rect 495102 672938 495134 673174
rect 494514 672854 495134 672938
rect 494514 672618 494546 672854
rect 494782 672618 494866 672854
rect 495102 672618 495134 672854
rect 494514 637174 495134 672618
rect 494514 636938 494546 637174
rect 494782 636938 494866 637174
rect 495102 636938 495134 637174
rect 494514 636854 495134 636938
rect 494514 636618 494546 636854
rect 494782 636618 494866 636854
rect 495102 636618 495134 636854
rect 494514 601174 495134 636618
rect 494514 600938 494546 601174
rect 494782 600938 494866 601174
rect 495102 600938 495134 601174
rect 494514 600854 495134 600938
rect 494514 600618 494546 600854
rect 494782 600618 494866 600854
rect 495102 600618 495134 600854
rect 494514 565174 495134 600618
rect 494514 564938 494546 565174
rect 494782 564938 494866 565174
rect 495102 564938 495134 565174
rect 494514 564854 495134 564938
rect 494514 564618 494546 564854
rect 494782 564618 494866 564854
rect 495102 564618 495134 564854
rect 494514 529174 495134 564618
rect 494514 528938 494546 529174
rect 494782 528938 494866 529174
rect 495102 528938 495134 529174
rect 494514 528854 495134 528938
rect 494514 528618 494546 528854
rect 494782 528618 494866 528854
rect 495102 528618 495134 528854
rect 494514 493174 495134 528618
rect 494514 492938 494546 493174
rect 494782 492938 494866 493174
rect 495102 492938 495134 493174
rect 494514 492854 495134 492938
rect 494514 492618 494546 492854
rect 494782 492618 494866 492854
rect 495102 492618 495134 492854
rect 494514 457174 495134 492618
rect 494514 456938 494546 457174
rect 494782 456938 494866 457174
rect 495102 456938 495134 457174
rect 494514 456854 495134 456938
rect 494514 456618 494546 456854
rect 494782 456618 494866 456854
rect 495102 456618 495134 456854
rect 494514 421174 495134 456618
rect 494514 420938 494546 421174
rect 494782 420938 494866 421174
rect 495102 420938 495134 421174
rect 494514 420854 495134 420938
rect 494514 420618 494546 420854
rect 494782 420618 494866 420854
rect 495102 420618 495134 420854
rect 494514 385174 495134 420618
rect 494514 384938 494546 385174
rect 494782 384938 494866 385174
rect 495102 384938 495134 385174
rect 494514 384854 495134 384938
rect 494514 384618 494546 384854
rect 494782 384618 494866 384854
rect 495102 384618 495134 384854
rect 494514 349174 495134 384618
rect 494514 348938 494546 349174
rect 494782 348938 494866 349174
rect 495102 348938 495134 349174
rect 494514 348854 495134 348938
rect 494514 348618 494546 348854
rect 494782 348618 494866 348854
rect 495102 348618 495134 348854
rect 494514 313174 495134 348618
rect 494514 312938 494546 313174
rect 494782 312938 494866 313174
rect 495102 312938 495134 313174
rect 494514 312854 495134 312938
rect 494514 312618 494546 312854
rect 494782 312618 494866 312854
rect 495102 312618 495134 312854
rect 494514 277174 495134 312618
rect 494514 276938 494546 277174
rect 494782 276938 494866 277174
rect 495102 276938 495134 277174
rect 494514 276854 495134 276938
rect 494514 276618 494546 276854
rect 494782 276618 494866 276854
rect 495102 276618 495134 276854
rect 494514 241174 495134 276618
rect 494514 240938 494546 241174
rect 494782 240938 494866 241174
rect 495102 240938 495134 241174
rect 494514 240854 495134 240938
rect 494514 240618 494546 240854
rect 494782 240618 494866 240854
rect 495102 240618 495134 240854
rect 494514 205174 495134 240618
rect 494514 204938 494546 205174
rect 494782 204938 494866 205174
rect 495102 204938 495134 205174
rect 494514 204854 495134 204938
rect 494514 204618 494546 204854
rect 494782 204618 494866 204854
rect 495102 204618 495134 204854
rect 494514 169174 495134 204618
rect 494514 168938 494546 169174
rect 494782 168938 494866 169174
rect 495102 168938 495134 169174
rect 494514 168854 495134 168938
rect 494514 168618 494546 168854
rect 494782 168618 494866 168854
rect 495102 168618 495134 168854
rect 494514 133174 495134 168618
rect 494514 132938 494546 133174
rect 494782 132938 494866 133174
rect 495102 132938 495134 133174
rect 494514 132854 495134 132938
rect 494514 132618 494546 132854
rect 494782 132618 494866 132854
rect 495102 132618 495134 132854
rect 494514 97174 495134 132618
rect 494514 96938 494546 97174
rect 494782 96938 494866 97174
rect 495102 96938 495134 97174
rect 494514 96854 495134 96938
rect 494514 96618 494546 96854
rect 494782 96618 494866 96854
rect 495102 96618 495134 96854
rect 494514 61174 495134 96618
rect 494514 60938 494546 61174
rect 494782 60938 494866 61174
rect 495102 60938 495134 61174
rect 494514 60854 495134 60938
rect 494514 60618 494546 60854
rect 494782 60618 494866 60854
rect 495102 60618 495134 60854
rect 494514 25174 495134 60618
rect 494514 24938 494546 25174
rect 494782 24938 494866 25174
rect 495102 24938 495134 25174
rect 494514 24854 495134 24938
rect 494514 24618 494546 24854
rect 494782 24618 494866 24854
rect 495102 24618 495134 24854
rect 494514 -3226 495134 24618
rect 494514 -3462 494546 -3226
rect 494782 -3462 494866 -3226
rect 495102 -3462 495134 -3226
rect 494514 -3546 495134 -3462
rect 494514 -3782 494546 -3546
rect 494782 -3782 494866 -3546
rect 495102 -3782 495134 -3546
rect 494514 -3814 495134 -3782
rect 498234 676894 498854 709082
rect 498234 676658 498266 676894
rect 498502 676658 498586 676894
rect 498822 676658 498854 676894
rect 498234 676574 498854 676658
rect 498234 676338 498266 676574
rect 498502 676338 498586 676574
rect 498822 676338 498854 676574
rect 498234 640894 498854 676338
rect 498234 640658 498266 640894
rect 498502 640658 498586 640894
rect 498822 640658 498854 640894
rect 498234 640574 498854 640658
rect 498234 640338 498266 640574
rect 498502 640338 498586 640574
rect 498822 640338 498854 640574
rect 498234 604894 498854 640338
rect 498234 604658 498266 604894
rect 498502 604658 498586 604894
rect 498822 604658 498854 604894
rect 498234 604574 498854 604658
rect 498234 604338 498266 604574
rect 498502 604338 498586 604574
rect 498822 604338 498854 604574
rect 498234 568894 498854 604338
rect 498234 568658 498266 568894
rect 498502 568658 498586 568894
rect 498822 568658 498854 568894
rect 498234 568574 498854 568658
rect 498234 568338 498266 568574
rect 498502 568338 498586 568574
rect 498822 568338 498854 568574
rect 498234 532894 498854 568338
rect 498234 532658 498266 532894
rect 498502 532658 498586 532894
rect 498822 532658 498854 532894
rect 498234 532574 498854 532658
rect 498234 532338 498266 532574
rect 498502 532338 498586 532574
rect 498822 532338 498854 532574
rect 498234 496894 498854 532338
rect 498234 496658 498266 496894
rect 498502 496658 498586 496894
rect 498822 496658 498854 496894
rect 498234 496574 498854 496658
rect 498234 496338 498266 496574
rect 498502 496338 498586 496574
rect 498822 496338 498854 496574
rect 498234 460894 498854 496338
rect 498234 460658 498266 460894
rect 498502 460658 498586 460894
rect 498822 460658 498854 460894
rect 498234 460574 498854 460658
rect 498234 460338 498266 460574
rect 498502 460338 498586 460574
rect 498822 460338 498854 460574
rect 498234 424894 498854 460338
rect 498234 424658 498266 424894
rect 498502 424658 498586 424894
rect 498822 424658 498854 424894
rect 498234 424574 498854 424658
rect 498234 424338 498266 424574
rect 498502 424338 498586 424574
rect 498822 424338 498854 424574
rect 498234 388894 498854 424338
rect 498234 388658 498266 388894
rect 498502 388658 498586 388894
rect 498822 388658 498854 388894
rect 498234 388574 498854 388658
rect 498234 388338 498266 388574
rect 498502 388338 498586 388574
rect 498822 388338 498854 388574
rect 498234 352894 498854 388338
rect 498234 352658 498266 352894
rect 498502 352658 498586 352894
rect 498822 352658 498854 352894
rect 498234 352574 498854 352658
rect 498234 352338 498266 352574
rect 498502 352338 498586 352574
rect 498822 352338 498854 352574
rect 498234 316894 498854 352338
rect 498234 316658 498266 316894
rect 498502 316658 498586 316894
rect 498822 316658 498854 316894
rect 498234 316574 498854 316658
rect 498234 316338 498266 316574
rect 498502 316338 498586 316574
rect 498822 316338 498854 316574
rect 498234 280894 498854 316338
rect 498234 280658 498266 280894
rect 498502 280658 498586 280894
rect 498822 280658 498854 280894
rect 498234 280574 498854 280658
rect 498234 280338 498266 280574
rect 498502 280338 498586 280574
rect 498822 280338 498854 280574
rect 498234 244894 498854 280338
rect 498234 244658 498266 244894
rect 498502 244658 498586 244894
rect 498822 244658 498854 244894
rect 498234 244574 498854 244658
rect 498234 244338 498266 244574
rect 498502 244338 498586 244574
rect 498822 244338 498854 244574
rect 498234 208894 498854 244338
rect 498234 208658 498266 208894
rect 498502 208658 498586 208894
rect 498822 208658 498854 208894
rect 498234 208574 498854 208658
rect 498234 208338 498266 208574
rect 498502 208338 498586 208574
rect 498822 208338 498854 208574
rect 498234 172894 498854 208338
rect 498234 172658 498266 172894
rect 498502 172658 498586 172894
rect 498822 172658 498854 172894
rect 498234 172574 498854 172658
rect 498234 172338 498266 172574
rect 498502 172338 498586 172574
rect 498822 172338 498854 172574
rect 498234 136894 498854 172338
rect 498234 136658 498266 136894
rect 498502 136658 498586 136894
rect 498822 136658 498854 136894
rect 498234 136574 498854 136658
rect 498234 136338 498266 136574
rect 498502 136338 498586 136574
rect 498822 136338 498854 136574
rect 498234 100894 498854 136338
rect 498234 100658 498266 100894
rect 498502 100658 498586 100894
rect 498822 100658 498854 100894
rect 498234 100574 498854 100658
rect 498234 100338 498266 100574
rect 498502 100338 498586 100574
rect 498822 100338 498854 100574
rect 498234 64894 498854 100338
rect 498234 64658 498266 64894
rect 498502 64658 498586 64894
rect 498822 64658 498854 64894
rect 498234 64574 498854 64658
rect 498234 64338 498266 64574
rect 498502 64338 498586 64574
rect 498822 64338 498854 64574
rect 498234 28894 498854 64338
rect 498234 28658 498266 28894
rect 498502 28658 498586 28894
rect 498822 28658 498854 28894
rect 498234 28574 498854 28658
rect 498234 28338 498266 28574
rect 498502 28338 498586 28574
rect 498822 28338 498854 28574
rect 498234 -5146 498854 28338
rect 500794 704838 501414 705830
rect 500794 704602 500826 704838
rect 501062 704602 501146 704838
rect 501382 704602 501414 704838
rect 500794 704518 501414 704602
rect 500794 704282 500826 704518
rect 501062 704282 501146 704518
rect 501382 704282 501414 704518
rect 500794 687454 501414 704282
rect 500794 687218 500826 687454
rect 501062 687218 501146 687454
rect 501382 687218 501414 687454
rect 500794 687134 501414 687218
rect 500794 686898 500826 687134
rect 501062 686898 501146 687134
rect 501382 686898 501414 687134
rect 500794 651454 501414 686898
rect 500794 651218 500826 651454
rect 501062 651218 501146 651454
rect 501382 651218 501414 651454
rect 500794 651134 501414 651218
rect 500794 650898 500826 651134
rect 501062 650898 501146 651134
rect 501382 650898 501414 651134
rect 500794 615454 501414 650898
rect 500794 615218 500826 615454
rect 501062 615218 501146 615454
rect 501382 615218 501414 615454
rect 500794 615134 501414 615218
rect 500794 614898 500826 615134
rect 501062 614898 501146 615134
rect 501382 614898 501414 615134
rect 500794 579454 501414 614898
rect 500794 579218 500826 579454
rect 501062 579218 501146 579454
rect 501382 579218 501414 579454
rect 500794 579134 501414 579218
rect 500794 578898 500826 579134
rect 501062 578898 501146 579134
rect 501382 578898 501414 579134
rect 500794 543454 501414 578898
rect 500794 543218 500826 543454
rect 501062 543218 501146 543454
rect 501382 543218 501414 543454
rect 500794 543134 501414 543218
rect 500794 542898 500826 543134
rect 501062 542898 501146 543134
rect 501382 542898 501414 543134
rect 500794 507454 501414 542898
rect 500794 507218 500826 507454
rect 501062 507218 501146 507454
rect 501382 507218 501414 507454
rect 500794 507134 501414 507218
rect 500794 506898 500826 507134
rect 501062 506898 501146 507134
rect 501382 506898 501414 507134
rect 500794 471454 501414 506898
rect 500794 471218 500826 471454
rect 501062 471218 501146 471454
rect 501382 471218 501414 471454
rect 500794 471134 501414 471218
rect 500794 470898 500826 471134
rect 501062 470898 501146 471134
rect 501382 470898 501414 471134
rect 500794 435454 501414 470898
rect 500794 435218 500826 435454
rect 501062 435218 501146 435454
rect 501382 435218 501414 435454
rect 500794 435134 501414 435218
rect 500794 434898 500826 435134
rect 501062 434898 501146 435134
rect 501382 434898 501414 435134
rect 500794 399454 501414 434898
rect 500794 399218 500826 399454
rect 501062 399218 501146 399454
rect 501382 399218 501414 399454
rect 500794 399134 501414 399218
rect 500794 398898 500826 399134
rect 501062 398898 501146 399134
rect 501382 398898 501414 399134
rect 500794 363454 501414 398898
rect 500794 363218 500826 363454
rect 501062 363218 501146 363454
rect 501382 363218 501414 363454
rect 500794 363134 501414 363218
rect 500794 362898 500826 363134
rect 501062 362898 501146 363134
rect 501382 362898 501414 363134
rect 500794 327454 501414 362898
rect 500794 327218 500826 327454
rect 501062 327218 501146 327454
rect 501382 327218 501414 327454
rect 500794 327134 501414 327218
rect 500794 326898 500826 327134
rect 501062 326898 501146 327134
rect 501382 326898 501414 327134
rect 500794 291454 501414 326898
rect 500794 291218 500826 291454
rect 501062 291218 501146 291454
rect 501382 291218 501414 291454
rect 500794 291134 501414 291218
rect 500794 290898 500826 291134
rect 501062 290898 501146 291134
rect 501382 290898 501414 291134
rect 500794 255454 501414 290898
rect 500794 255218 500826 255454
rect 501062 255218 501146 255454
rect 501382 255218 501414 255454
rect 500794 255134 501414 255218
rect 500794 254898 500826 255134
rect 501062 254898 501146 255134
rect 501382 254898 501414 255134
rect 500794 219454 501414 254898
rect 500794 219218 500826 219454
rect 501062 219218 501146 219454
rect 501382 219218 501414 219454
rect 500794 219134 501414 219218
rect 500794 218898 500826 219134
rect 501062 218898 501146 219134
rect 501382 218898 501414 219134
rect 500794 183454 501414 218898
rect 500794 183218 500826 183454
rect 501062 183218 501146 183454
rect 501382 183218 501414 183454
rect 500794 183134 501414 183218
rect 500794 182898 500826 183134
rect 501062 182898 501146 183134
rect 501382 182898 501414 183134
rect 500794 147454 501414 182898
rect 500794 147218 500826 147454
rect 501062 147218 501146 147454
rect 501382 147218 501414 147454
rect 500794 147134 501414 147218
rect 500794 146898 500826 147134
rect 501062 146898 501146 147134
rect 501382 146898 501414 147134
rect 500794 111454 501414 146898
rect 500794 111218 500826 111454
rect 501062 111218 501146 111454
rect 501382 111218 501414 111454
rect 500794 111134 501414 111218
rect 500794 110898 500826 111134
rect 501062 110898 501146 111134
rect 501382 110898 501414 111134
rect 500794 75454 501414 110898
rect 500794 75218 500826 75454
rect 501062 75218 501146 75454
rect 501382 75218 501414 75454
rect 500794 75134 501414 75218
rect 500794 74898 500826 75134
rect 501062 74898 501146 75134
rect 501382 74898 501414 75134
rect 500794 39454 501414 74898
rect 500794 39218 500826 39454
rect 501062 39218 501146 39454
rect 501382 39218 501414 39454
rect 500794 39134 501414 39218
rect 500794 38898 500826 39134
rect 501062 38898 501146 39134
rect 501382 38898 501414 39134
rect 500794 3454 501414 38898
rect 500794 3218 500826 3454
rect 501062 3218 501146 3454
rect 501382 3218 501414 3454
rect 500794 3134 501414 3218
rect 500794 2898 500826 3134
rect 501062 2898 501146 3134
rect 501382 2898 501414 3134
rect 500794 -346 501414 2898
rect 500794 -582 500826 -346
rect 501062 -582 501146 -346
rect 501382 -582 501414 -346
rect 500794 -666 501414 -582
rect 500794 -902 500826 -666
rect 501062 -902 501146 -666
rect 501382 -902 501414 -666
rect 500794 -1894 501414 -902
rect 501954 680614 502574 711002
rect 511954 710598 512574 711590
rect 511954 710362 511986 710598
rect 512222 710362 512306 710598
rect 512542 710362 512574 710598
rect 511954 710278 512574 710362
rect 511954 710042 511986 710278
rect 512222 710042 512306 710278
rect 512542 710042 512574 710278
rect 508234 708678 508854 709670
rect 508234 708442 508266 708678
rect 508502 708442 508586 708678
rect 508822 708442 508854 708678
rect 508234 708358 508854 708442
rect 508234 708122 508266 708358
rect 508502 708122 508586 708358
rect 508822 708122 508854 708358
rect 501954 680378 501986 680614
rect 502222 680378 502306 680614
rect 502542 680378 502574 680614
rect 501954 680294 502574 680378
rect 501954 680058 501986 680294
rect 502222 680058 502306 680294
rect 502542 680058 502574 680294
rect 501954 644614 502574 680058
rect 501954 644378 501986 644614
rect 502222 644378 502306 644614
rect 502542 644378 502574 644614
rect 501954 644294 502574 644378
rect 501954 644058 501986 644294
rect 502222 644058 502306 644294
rect 502542 644058 502574 644294
rect 501954 608614 502574 644058
rect 501954 608378 501986 608614
rect 502222 608378 502306 608614
rect 502542 608378 502574 608614
rect 501954 608294 502574 608378
rect 501954 608058 501986 608294
rect 502222 608058 502306 608294
rect 502542 608058 502574 608294
rect 501954 572614 502574 608058
rect 501954 572378 501986 572614
rect 502222 572378 502306 572614
rect 502542 572378 502574 572614
rect 501954 572294 502574 572378
rect 501954 572058 501986 572294
rect 502222 572058 502306 572294
rect 502542 572058 502574 572294
rect 501954 536614 502574 572058
rect 501954 536378 501986 536614
rect 502222 536378 502306 536614
rect 502542 536378 502574 536614
rect 501954 536294 502574 536378
rect 501954 536058 501986 536294
rect 502222 536058 502306 536294
rect 502542 536058 502574 536294
rect 501954 500614 502574 536058
rect 501954 500378 501986 500614
rect 502222 500378 502306 500614
rect 502542 500378 502574 500614
rect 501954 500294 502574 500378
rect 501954 500058 501986 500294
rect 502222 500058 502306 500294
rect 502542 500058 502574 500294
rect 501954 464614 502574 500058
rect 501954 464378 501986 464614
rect 502222 464378 502306 464614
rect 502542 464378 502574 464614
rect 501954 464294 502574 464378
rect 501954 464058 501986 464294
rect 502222 464058 502306 464294
rect 502542 464058 502574 464294
rect 501954 428614 502574 464058
rect 501954 428378 501986 428614
rect 502222 428378 502306 428614
rect 502542 428378 502574 428614
rect 501954 428294 502574 428378
rect 501954 428058 501986 428294
rect 502222 428058 502306 428294
rect 502542 428058 502574 428294
rect 501954 392614 502574 428058
rect 501954 392378 501986 392614
rect 502222 392378 502306 392614
rect 502542 392378 502574 392614
rect 501954 392294 502574 392378
rect 501954 392058 501986 392294
rect 502222 392058 502306 392294
rect 502542 392058 502574 392294
rect 501954 356614 502574 392058
rect 501954 356378 501986 356614
rect 502222 356378 502306 356614
rect 502542 356378 502574 356614
rect 501954 356294 502574 356378
rect 501954 356058 501986 356294
rect 502222 356058 502306 356294
rect 502542 356058 502574 356294
rect 501954 320614 502574 356058
rect 501954 320378 501986 320614
rect 502222 320378 502306 320614
rect 502542 320378 502574 320614
rect 501954 320294 502574 320378
rect 501954 320058 501986 320294
rect 502222 320058 502306 320294
rect 502542 320058 502574 320294
rect 501954 284614 502574 320058
rect 501954 284378 501986 284614
rect 502222 284378 502306 284614
rect 502542 284378 502574 284614
rect 501954 284294 502574 284378
rect 501954 284058 501986 284294
rect 502222 284058 502306 284294
rect 502542 284058 502574 284294
rect 501954 248614 502574 284058
rect 501954 248378 501986 248614
rect 502222 248378 502306 248614
rect 502542 248378 502574 248614
rect 501954 248294 502574 248378
rect 501954 248058 501986 248294
rect 502222 248058 502306 248294
rect 502542 248058 502574 248294
rect 501954 212614 502574 248058
rect 501954 212378 501986 212614
rect 502222 212378 502306 212614
rect 502542 212378 502574 212614
rect 501954 212294 502574 212378
rect 501954 212058 501986 212294
rect 502222 212058 502306 212294
rect 502542 212058 502574 212294
rect 501954 176614 502574 212058
rect 501954 176378 501986 176614
rect 502222 176378 502306 176614
rect 502542 176378 502574 176614
rect 501954 176294 502574 176378
rect 501954 176058 501986 176294
rect 502222 176058 502306 176294
rect 502542 176058 502574 176294
rect 501954 140614 502574 176058
rect 501954 140378 501986 140614
rect 502222 140378 502306 140614
rect 502542 140378 502574 140614
rect 501954 140294 502574 140378
rect 501954 140058 501986 140294
rect 502222 140058 502306 140294
rect 502542 140058 502574 140294
rect 501954 104614 502574 140058
rect 501954 104378 501986 104614
rect 502222 104378 502306 104614
rect 502542 104378 502574 104614
rect 501954 104294 502574 104378
rect 501954 104058 501986 104294
rect 502222 104058 502306 104294
rect 502542 104058 502574 104294
rect 501954 68614 502574 104058
rect 501954 68378 501986 68614
rect 502222 68378 502306 68614
rect 502542 68378 502574 68614
rect 501954 68294 502574 68378
rect 501954 68058 501986 68294
rect 502222 68058 502306 68294
rect 502542 68058 502574 68294
rect 501954 32614 502574 68058
rect 501954 32378 501986 32614
rect 502222 32378 502306 32614
rect 502542 32378 502574 32614
rect 501954 32294 502574 32378
rect 501954 32058 501986 32294
rect 502222 32058 502306 32294
rect 502542 32058 502574 32294
rect 498234 -5382 498266 -5146
rect 498502 -5382 498586 -5146
rect 498822 -5382 498854 -5146
rect 498234 -5466 498854 -5382
rect 498234 -5702 498266 -5466
rect 498502 -5702 498586 -5466
rect 498822 -5702 498854 -5466
rect 498234 -5734 498854 -5702
rect 491954 -6342 491986 -6106
rect 492222 -6342 492306 -6106
rect 492542 -6342 492574 -6106
rect 491954 -6426 492574 -6342
rect 491954 -6662 491986 -6426
rect 492222 -6662 492306 -6426
rect 492542 -6662 492574 -6426
rect 491954 -7654 492574 -6662
rect 501954 -7066 502574 32058
rect 504514 706758 505134 707750
rect 504514 706522 504546 706758
rect 504782 706522 504866 706758
rect 505102 706522 505134 706758
rect 504514 706438 505134 706522
rect 504514 706202 504546 706438
rect 504782 706202 504866 706438
rect 505102 706202 505134 706438
rect 504514 691174 505134 706202
rect 504514 690938 504546 691174
rect 504782 690938 504866 691174
rect 505102 690938 505134 691174
rect 504514 690854 505134 690938
rect 504514 690618 504546 690854
rect 504782 690618 504866 690854
rect 505102 690618 505134 690854
rect 504514 655174 505134 690618
rect 504514 654938 504546 655174
rect 504782 654938 504866 655174
rect 505102 654938 505134 655174
rect 504514 654854 505134 654938
rect 504514 654618 504546 654854
rect 504782 654618 504866 654854
rect 505102 654618 505134 654854
rect 504514 619174 505134 654618
rect 504514 618938 504546 619174
rect 504782 618938 504866 619174
rect 505102 618938 505134 619174
rect 504514 618854 505134 618938
rect 504514 618618 504546 618854
rect 504782 618618 504866 618854
rect 505102 618618 505134 618854
rect 504514 583174 505134 618618
rect 504514 582938 504546 583174
rect 504782 582938 504866 583174
rect 505102 582938 505134 583174
rect 504514 582854 505134 582938
rect 504514 582618 504546 582854
rect 504782 582618 504866 582854
rect 505102 582618 505134 582854
rect 504514 547174 505134 582618
rect 504514 546938 504546 547174
rect 504782 546938 504866 547174
rect 505102 546938 505134 547174
rect 504514 546854 505134 546938
rect 504514 546618 504546 546854
rect 504782 546618 504866 546854
rect 505102 546618 505134 546854
rect 504514 511174 505134 546618
rect 504514 510938 504546 511174
rect 504782 510938 504866 511174
rect 505102 510938 505134 511174
rect 504514 510854 505134 510938
rect 504514 510618 504546 510854
rect 504782 510618 504866 510854
rect 505102 510618 505134 510854
rect 504514 475174 505134 510618
rect 504514 474938 504546 475174
rect 504782 474938 504866 475174
rect 505102 474938 505134 475174
rect 504514 474854 505134 474938
rect 504514 474618 504546 474854
rect 504782 474618 504866 474854
rect 505102 474618 505134 474854
rect 504514 439174 505134 474618
rect 504514 438938 504546 439174
rect 504782 438938 504866 439174
rect 505102 438938 505134 439174
rect 504514 438854 505134 438938
rect 504514 438618 504546 438854
rect 504782 438618 504866 438854
rect 505102 438618 505134 438854
rect 504514 403174 505134 438618
rect 504514 402938 504546 403174
rect 504782 402938 504866 403174
rect 505102 402938 505134 403174
rect 504514 402854 505134 402938
rect 504514 402618 504546 402854
rect 504782 402618 504866 402854
rect 505102 402618 505134 402854
rect 504514 367174 505134 402618
rect 504514 366938 504546 367174
rect 504782 366938 504866 367174
rect 505102 366938 505134 367174
rect 504514 366854 505134 366938
rect 504514 366618 504546 366854
rect 504782 366618 504866 366854
rect 505102 366618 505134 366854
rect 504514 331174 505134 366618
rect 504514 330938 504546 331174
rect 504782 330938 504866 331174
rect 505102 330938 505134 331174
rect 504514 330854 505134 330938
rect 504514 330618 504546 330854
rect 504782 330618 504866 330854
rect 505102 330618 505134 330854
rect 504514 295174 505134 330618
rect 504514 294938 504546 295174
rect 504782 294938 504866 295174
rect 505102 294938 505134 295174
rect 504514 294854 505134 294938
rect 504514 294618 504546 294854
rect 504782 294618 504866 294854
rect 505102 294618 505134 294854
rect 504514 259174 505134 294618
rect 504514 258938 504546 259174
rect 504782 258938 504866 259174
rect 505102 258938 505134 259174
rect 504514 258854 505134 258938
rect 504514 258618 504546 258854
rect 504782 258618 504866 258854
rect 505102 258618 505134 258854
rect 504514 223174 505134 258618
rect 504514 222938 504546 223174
rect 504782 222938 504866 223174
rect 505102 222938 505134 223174
rect 504514 222854 505134 222938
rect 504514 222618 504546 222854
rect 504782 222618 504866 222854
rect 505102 222618 505134 222854
rect 504514 187174 505134 222618
rect 504514 186938 504546 187174
rect 504782 186938 504866 187174
rect 505102 186938 505134 187174
rect 504514 186854 505134 186938
rect 504514 186618 504546 186854
rect 504782 186618 504866 186854
rect 505102 186618 505134 186854
rect 504514 151174 505134 186618
rect 504514 150938 504546 151174
rect 504782 150938 504866 151174
rect 505102 150938 505134 151174
rect 504514 150854 505134 150938
rect 504514 150618 504546 150854
rect 504782 150618 504866 150854
rect 505102 150618 505134 150854
rect 504514 115174 505134 150618
rect 504514 114938 504546 115174
rect 504782 114938 504866 115174
rect 505102 114938 505134 115174
rect 504514 114854 505134 114938
rect 504514 114618 504546 114854
rect 504782 114618 504866 114854
rect 505102 114618 505134 114854
rect 504514 79174 505134 114618
rect 504514 78938 504546 79174
rect 504782 78938 504866 79174
rect 505102 78938 505134 79174
rect 504514 78854 505134 78938
rect 504514 78618 504546 78854
rect 504782 78618 504866 78854
rect 505102 78618 505134 78854
rect 504514 43174 505134 78618
rect 504514 42938 504546 43174
rect 504782 42938 504866 43174
rect 505102 42938 505134 43174
rect 504514 42854 505134 42938
rect 504514 42618 504546 42854
rect 504782 42618 504866 42854
rect 505102 42618 505134 42854
rect 504514 7174 505134 42618
rect 504514 6938 504546 7174
rect 504782 6938 504866 7174
rect 505102 6938 505134 7174
rect 504514 6854 505134 6938
rect 504514 6618 504546 6854
rect 504782 6618 504866 6854
rect 505102 6618 505134 6854
rect 504514 -2266 505134 6618
rect 504514 -2502 504546 -2266
rect 504782 -2502 504866 -2266
rect 505102 -2502 505134 -2266
rect 504514 -2586 505134 -2502
rect 504514 -2822 504546 -2586
rect 504782 -2822 504866 -2586
rect 505102 -2822 505134 -2586
rect 504514 -3814 505134 -2822
rect 508234 694894 508854 708122
rect 508234 694658 508266 694894
rect 508502 694658 508586 694894
rect 508822 694658 508854 694894
rect 508234 694574 508854 694658
rect 508234 694338 508266 694574
rect 508502 694338 508586 694574
rect 508822 694338 508854 694574
rect 508234 658894 508854 694338
rect 508234 658658 508266 658894
rect 508502 658658 508586 658894
rect 508822 658658 508854 658894
rect 508234 658574 508854 658658
rect 508234 658338 508266 658574
rect 508502 658338 508586 658574
rect 508822 658338 508854 658574
rect 508234 622894 508854 658338
rect 508234 622658 508266 622894
rect 508502 622658 508586 622894
rect 508822 622658 508854 622894
rect 508234 622574 508854 622658
rect 508234 622338 508266 622574
rect 508502 622338 508586 622574
rect 508822 622338 508854 622574
rect 508234 586894 508854 622338
rect 508234 586658 508266 586894
rect 508502 586658 508586 586894
rect 508822 586658 508854 586894
rect 508234 586574 508854 586658
rect 508234 586338 508266 586574
rect 508502 586338 508586 586574
rect 508822 586338 508854 586574
rect 508234 550894 508854 586338
rect 508234 550658 508266 550894
rect 508502 550658 508586 550894
rect 508822 550658 508854 550894
rect 508234 550574 508854 550658
rect 508234 550338 508266 550574
rect 508502 550338 508586 550574
rect 508822 550338 508854 550574
rect 508234 514894 508854 550338
rect 508234 514658 508266 514894
rect 508502 514658 508586 514894
rect 508822 514658 508854 514894
rect 508234 514574 508854 514658
rect 508234 514338 508266 514574
rect 508502 514338 508586 514574
rect 508822 514338 508854 514574
rect 508234 478894 508854 514338
rect 508234 478658 508266 478894
rect 508502 478658 508586 478894
rect 508822 478658 508854 478894
rect 508234 478574 508854 478658
rect 508234 478338 508266 478574
rect 508502 478338 508586 478574
rect 508822 478338 508854 478574
rect 508234 442894 508854 478338
rect 508234 442658 508266 442894
rect 508502 442658 508586 442894
rect 508822 442658 508854 442894
rect 508234 442574 508854 442658
rect 508234 442338 508266 442574
rect 508502 442338 508586 442574
rect 508822 442338 508854 442574
rect 508234 406894 508854 442338
rect 508234 406658 508266 406894
rect 508502 406658 508586 406894
rect 508822 406658 508854 406894
rect 508234 406574 508854 406658
rect 508234 406338 508266 406574
rect 508502 406338 508586 406574
rect 508822 406338 508854 406574
rect 508234 370894 508854 406338
rect 508234 370658 508266 370894
rect 508502 370658 508586 370894
rect 508822 370658 508854 370894
rect 508234 370574 508854 370658
rect 508234 370338 508266 370574
rect 508502 370338 508586 370574
rect 508822 370338 508854 370574
rect 508234 334894 508854 370338
rect 508234 334658 508266 334894
rect 508502 334658 508586 334894
rect 508822 334658 508854 334894
rect 508234 334574 508854 334658
rect 508234 334338 508266 334574
rect 508502 334338 508586 334574
rect 508822 334338 508854 334574
rect 508234 298894 508854 334338
rect 508234 298658 508266 298894
rect 508502 298658 508586 298894
rect 508822 298658 508854 298894
rect 508234 298574 508854 298658
rect 508234 298338 508266 298574
rect 508502 298338 508586 298574
rect 508822 298338 508854 298574
rect 508234 262894 508854 298338
rect 508234 262658 508266 262894
rect 508502 262658 508586 262894
rect 508822 262658 508854 262894
rect 508234 262574 508854 262658
rect 508234 262338 508266 262574
rect 508502 262338 508586 262574
rect 508822 262338 508854 262574
rect 508234 226894 508854 262338
rect 508234 226658 508266 226894
rect 508502 226658 508586 226894
rect 508822 226658 508854 226894
rect 508234 226574 508854 226658
rect 508234 226338 508266 226574
rect 508502 226338 508586 226574
rect 508822 226338 508854 226574
rect 508234 190894 508854 226338
rect 508234 190658 508266 190894
rect 508502 190658 508586 190894
rect 508822 190658 508854 190894
rect 508234 190574 508854 190658
rect 508234 190338 508266 190574
rect 508502 190338 508586 190574
rect 508822 190338 508854 190574
rect 508234 154894 508854 190338
rect 508234 154658 508266 154894
rect 508502 154658 508586 154894
rect 508822 154658 508854 154894
rect 508234 154574 508854 154658
rect 508234 154338 508266 154574
rect 508502 154338 508586 154574
rect 508822 154338 508854 154574
rect 508234 118894 508854 154338
rect 508234 118658 508266 118894
rect 508502 118658 508586 118894
rect 508822 118658 508854 118894
rect 508234 118574 508854 118658
rect 508234 118338 508266 118574
rect 508502 118338 508586 118574
rect 508822 118338 508854 118574
rect 508234 82894 508854 118338
rect 508234 82658 508266 82894
rect 508502 82658 508586 82894
rect 508822 82658 508854 82894
rect 508234 82574 508854 82658
rect 508234 82338 508266 82574
rect 508502 82338 508586 82574
rect 508822 82338 508854 82574
rect 508234 46894 508854 82338
rect 508234 46658 508266 46894
rect 508502 46658 508586 46894
rect 508822 46658 508854 46894
rect 508234 46574 508854 46658
rect 508234 46338 508266 46574
rect 508502 46338 508586 46574
rect 508822 46338 508854 46574
rect 508234 10894 508854 46338
rect 508234 10658 508266 10894
rect 508502 10658 508586 10894
rect 508822 10658 508854 10894
rect 508234 10574 508854 10658
rect 508234 10338 508266 10574
rect 508502 10338 508586 10574
rect 508822 10338 508854 10574
rect 508234 -4186 508854 10338
rect 510794 705798 511414 705830
rect 510794 705562 510826 705798
rect 511062 705562 511146 705798
rect 511382 705562 511414 705798
rect 510794 705478 511414 705562
rect 510794 705242 510826 705478
rect 511062 705242 511146 705478
rect 511382 705242 511414 705478
rect 510794 669454 511414 705242
rect 510794 669218 510826 669454
rect 511062 669218 511146 669454
rect 511382 669218 511414 669454
rect 510794 669134 511414 669218
rect 510794 668898 510826 669134
rect 511062 668898 511146 669134
rect 511382 668898 511414 669134
rect 510794 633454 511414 668898
rect 510794 633218 510826 633454
rect 511062 633218 511146 633454
rect 511382 633218 511414 633454
rect 510794 633134 511414 633218
rect 510794 632898 510826 633134
rect 511062 632898 511146 633134
rect 511382 632898 511414 633134
rect 510794 597454 511414 632898
rect 510794 597218 510826 597454
rect 511062 597218 511146 597454
rect 511382 597218 511414 597454
rect 510794 597134 511414 597218
rect 510794 596898 510826 597134
rect 511062 596898 511146 597134
rect 511382 596898 511414 597134
rect 510794 561454 511414 596898
rect 510794 561218 510826 561454
rect 511062 561218 511146 561454
rect 511382 561218 511414 561454
rect 510794 561134 511414 561218
rect 510794 560898 510826 561134
rect 511062 560898 511146 561134
rect 511382 560898 511414 561134
rect 510794 525454 511414 560898
rect 510794 525218 510826 525454
rect 511062 525218 511146 525454
rect 511382 525218 511414 525454
rect 510794 525134 511414 525218
rect 510794 524898 510826 525134
rect 511062 524898 511146 525134
rect 511382 524898 511414 525134
rect 510794 489454 511414 524898
rect 510794 489218 510826 489454
rect 511062 489218 511146 489454
rect 511382 489218 511414 489454
rect 510794 489134 511414 489218
rect 510794 488898 510826 489134
rect 511062 488898 511146 489134
rect 511382 488898 511414 489134
rect 510794 453454 511414 488898
rect 510794 453218 510826 453454
rect 511062 453218 511146 453454
rect 511382 453218 511414 453454
rect 510794 453134 511414 453218
rect 510794 452898 510826 453134
rect 511062 452898 511146 453134
rect 511382 452898 511414 453134
rect 510794 417454 511414 452898
rect 510794 417218 510826 417454
rect 511062 417218 511146 417454
rect 511382 417218 511414 417454
rect 510794 417134 511414 417218
rect 510794 416898 510826 417134
rect 511062 416898 511146 417134
rect 511382 416898 511414 417134
rect 510794 381454 511414 416898
rect 510794 381218 510826 381454
rect 511062 381218 511146 381454
rect 511382 381218 511414 381454
rect 510794 381134 511414 381218
rect 510794 380898 510826 381134
rect 511062 380898 511146 381134
rect 511382 380898 511414 381134
rect 510794 345454 511414 380898
rect 510794 345218 510826 345454
rect 511062 345218 511146 345454
rect 511382 345218 511414 345454
rect 510794 345134 511414 345218
rect 510794 344898 510826 345134
rect 511062 344898 511146 345134
rect 511382 344898 511414 345134
rect 510794 309454 511414 344898
rect 510794 309218 510826 309454
rect 511062 309218 511146 309454
rect 511382 309218 511414 309454
rect 510794 309134 511414 309218
rect 510794 308898 510826 309134
rect 511062 308898 511146 309134
rect 511382 308898 511414 309134
rect 510794 273454 511414 308898
rect 510794 273218 510826 273454
rect 511062 273218 511146 273454
rect 511382 273218 511414 273454
rect 510794 273134 511414 273218
rect 510794 272898 510826 273134
rect 511062 272898 511146 273134
rect 511382 272898 511414 273134
rect 510794 237454 511414 272898
rect 510794 237218 510826 237454
rect 511062 237218 511146 237454
rect 511382 237218 511414 237454
rect 510794 237134 511414 237218
rect 510794 236898 510826 237134
rect 511062 236898 511146 237134
rect 511382 236898 511414 237134
rect 510794 201454 511414 236898
rect 510794 201218 510826 201454
rect 511062 201218 511146 201454
rect 511382 201218 511414 201454
rect 510794 201134 511414 201218
rect 510794 200898 510826 201134
rect 511062 200898 511146 201134
rect 511382 200898 511414 201134
rect 510794 165454 511414 200898
rect 510794 165218 510826 165454
rect 511062 165218 511146 165454
rect 511382 165218 511414 165454
rect 510794 165134 511414 165218
rect 510794 164898 510826 165134
rect 511062 164898 511146 165134
rect 511382 164898 511414 165134
rect 510794 129454 511414 164898
rect 510794 129218 510826 129454
rect 511062 129218 511146 129454
rect 511382 129218 511414 129454
rect 510794 129134 511414 129218
rect 510794 128898 510826 129134
rect 511062 128898 511146 129134
rect 511382 128898 511414 129134
rect 510794 93454 511414 128898
rect 510794 93218 510826 93454
rect 511062 93218 511146 93454
rect 511382 93218 511414 93454
rect 510794 93134 511414 93218
rect 510794 92898 510826 93134
rect 511062 92898 511146 93134
rect 511382 92898 511414 93134
rect 510794 57454 511414 92898
rect 510794 57218 510826 57454
rect 511062 57218 511146 57454
rect 511382 57218 511414 57454
rect 510794 57134 511414 57218
rect 510794 56898 510826 57134
rect 511062 56898 511146 57134
rect 511382 56898 511414 57134
rect 510794 21454 511414 56898
rect 510794 21218 510826 21454
rect 511062 21218 511146 21454
rect 511382 21218 511414 21454
rect 510794 21134 511414 21218
rect 510794 20898 510826 21134
rect 511062 20898 511146 21134
rect 511382 20898 511414 21134
rect 510794 -1306 511414 20898
rect 510794 -1542 510826 -1306
rect 511062 -1542 511146 -1306
rect 511382 -1542 511414 -1306
rect 510794 -1626 511414 -1542
rect 510794 -1862 510826 -1626
rect 511062 -1862 511146 -1626
rect 511382 -1862 511414 -1626
rect 510794 -1894 511414 -1862
rect 511954 698614 512574 710042
rect 521954 711558 522574 711590
rect 521954 711322 521986 711558
rect 522222 711322 522306 711558
rect 522542 711322 522574 711558
rect 521954 711238 522574 711322
rect 521954 711002 521986 711238
rect 522222 711002 522306 711238
rect 522542 711002 522574 711238
rect 518234 709638 518854 709670
rect 518234 709402 518266 709638
rect 518502 709402 518586 709638
rect 518822 709402 518854 709638
rect 518234 709318 518854 709402
rect 518234 709082 518266 709318
rect 518502 709082 518586 709318
rect 518822 709082 518854 709318
rect 511954 698378 511986 698614
rect 512222 698378 512306 698614
rect 512542 698378 512574 698614
rect 511954 698294 512574 698378
rect 511954 698058 511986 698294
rect 512222 698058 512306 698294
rect 512542 698058 512574 698294
rect 511954 662614 512574 698058
rect 511954 662378 511986 662614
rect 512222 662378 512306 662614
rect 512542 662378 512574 662614
rect 511954 662294 512574 662378
rect 511954 662058 511986 662294
rect 512222 662058 512306 662294
rect 512542 662058 512574 662294
rect 511954 626614 512574 662058
rect 511954 626378 511986 626614
rect 512222 626378 512306 626614
rect 512542 626378 512574 626614
rect 511954 626294 512574 626378
rect 511954 626058 511986 626294
rect 512222 626058 512306 626294
rect 512542 626058 512574 626294
rect 511954 590614 512574 626058
rect 511954 590378 511986 590614
rect 512222 590378 512306 590614
rect 512542 590378 512574 590614
rect 511954 590294 512574 590378
rect 511954 590058 511986 590294
rect 512222 590058 512306 590294
rect 512542 590058 512574 590294
rect 511954 554614 512574 590058
rect 511954 554378 511986 554614
rect 512222 554378 512306 554614
rect 512542 554378 512574 554614
rect 511954 554294 512574 554378
rect 511954 554058 511986 554294
rect 512222 554058 512306 554294
rect 512542 554058 512574 554294
rect 511954 518614 512574 554058
rect 511954 518378 511986 518614
rect 512222 518378 512306 518614
rect 512542 518378 512574 518614
rect 511954 518294 512574 518378
rect 511954 518058 511986 518294
rect 512222 518058 512306 518294
rect 512542 518058 512574 518294
rect 511954 482614 512574 518058
rect 511954 482378 511986 482614
rect 512222 482378 512306 482614
rect 512542 482378 512574 482614
rect 511954 482294 512574 482378
rect 511954 482058 511986 482294
rect 512222 482058 512306 482294
rect 512542 482058 512574 482294
rect 511954 446614 512574 482058
rect 511954 446378 511986 446614
rect 512222 446378 512306 446614
rect 512542 446378 512574 446614
rect 511954 446294 512574 446378
rect 511954 446058 511986 446294
rect 512222 446058 512306 446294
rect 512542 446058 512574 446294
rect 511954 410614 512574 446058
rect 511954 410378 511986 410614
rect 512222 410378 512306 410614
rect 512542 410378 512574 410614
rect 511954 410294 512574 410378
rect 511954 410058 511986 410294
rect 512222 410058 512306 410294
rect 512542 410058 512574 410294
rect 511954 374614 512574 410058
rect 511954 374378 511986 374614
rect 512222 374378 512306 374614
rect 512542 374378 512574 374614
rect 511954 374294 512574 374378
rect 511954 374058 511986 374294
rect 512222 374058 512306 374294
rect 512542 374058 512574 374294
rect 511954 338614 512574 374058
rect 511954 338378 511986 338614
rect 512222 338378 512306 338614
rect 512542 338378 512574 338614
rect 511954 338294 512574 338378
rect 511954 338058 511986 338294
rect 512222 338058 512306 338294
rect 512542 338058 512574 338294
rect 511954 302614 512574 338058
rect 511954 302378 511986 302614
rect 512222 302378 512306 302614
rect 512542 302378 512574 302614
rect 511954 302294 512574 302378
rect 511954 302058 511986 302294
rect 512222 302058 512306 302294
rect 512542 302058 512574 302294
rect 511954 266614 512574 302058
rect 511954 266378 511986 266614
rect 512222 266378 512306 266614
rect 512542 266378 512574 266614
rect 511954 266294 512574 266378
rect 511954 266058 511986 266294
rect 512222 266058 512306 266294
rect 512542 266058 512574 266294
rect 511954 230614 512574 266058
rect 511954 230378 511986 230614
rect 512222 230378 512306 230614
rect 512542 230378 512574 230614
rect 511954 230294 512574 230378
rect 511954 230058 511986 230294
rect 512222 230058 512306 230294
rect 512542 230058 512574 230294
rect 511954 194614 512574 230058
rect 511954 194378 511986 194614
rect 512222 194378 512306 194614
rect 512542 194378 512574 194614
rect 511954 194294 512574 194378
rect 511954 194058 511986 194294
rect 512222 194058 512306 194294
rect 512542 194058 512574 194294
rect 511954 158614 512574 194058
rect 511954 158378 511986 158614
rect 512222 158378 512306 158614
rect 512542 158378 512574 158614
rect 511954 158294 512574 158378
rect 511954 158058 511986 158294
rect 512222 158058 512306 158294
rect 512542 158058 512574 158294
rect 511954 122614 512574 158058
rect 511954 122378 511986 122614
rect 512222 122378 512306 122614
rect 512542 122378 512574 122614
rect 511954 122294 512574 122378
rect 511954 122058 511986 122294
rect 512222 122058 512306 122294
rect 512542 122058 512574 122294
rect 511954 86614 512574 122058
rect 511954 86378 511986 86614
rect 512222 86378 512306 86614
rect 512542 86378 512574 86614
rect 511954 86294 512574 86378
rect 511954 86058 511986 86294
rect 512222 86058 512306 86294
rect 512542 86058 512574 86294
rect 511954 50614 512574 86058
rect 511954 50378 511986 50614
rect 512222 50378 512306 50614
rect 512542 50378 512574 50614
rect 511954 50294 512574 50378
rect 511954 50058 511986 50294
rect 512222 50058 512306 50294
rect 512542 50058 512574 50294
rect 511954 14614 512574 50058
rect 511954 14378 511986 14614
rect 512222 14378 512306 14614
rect 512542 14378 512574 14614
rect 511954 14294 512574 14378
rect 511954 14058 511986 14294
rect 512222 14058 512306 14294
rect 512542 14058 512574 14294
rect 508234 -4422 508266 -4186
rect 508502 -4422 508586 -4186
rect 508822 -4422 508854 -4186
rect 508234 -4506 508854 -4422
rect 508234 -4742 508266 -4506
rect 508502 -4742 508586 -4506
rect 508822 -4742 508854 -4506
rect 508234 -5734 508854 -4742
rect 501954 -7302 501986 -7066
rect 502222 -7302 502306 -7066
rect 502542 -7302 502574 -7066
rect 501954 -7386 502574 -7302
rect 501954 -7622 501986 -7386
rect 502222 -7622 502306 -7386
rect 502542 -7622 502574 -7386
rect 501954 -7654 502574 -7622
rect 511954 -6106 512574 14058
rect 514514 707718 515134 707750
rect 514514 707482 514546 707718
rect 514782 707482 514866 707718
rect 515102 707482 515134 707718
rect 514514 707398 515134 707482
rect 514514 707162 514546 707398
rect 514782 707162 514866 707398
rect 515102 707162 515134 707398
rect 514514 673174 515134 707162
rect 514514 672938 514546 673174
rect 514782 672938 514866 673174
rect 515102 672938 515134 673174
rect 514514 672854 515134 672938
rect 514514 672618 514546 672854
rect 514782 672618 514866 672854
rect 515102 672618 515134 672854
rect 514514 637174 515134 672618
rect 514514 636938 514546 637174
rect 514782 636938 514866 637174
rect 515102 636938 515134 637174
rect 514514 636854 515134 636938
rect 514514 636618 514546 636854
rect 514782 636618 514866 636854
rect 515102 636618 515134 636854
rect 514514 601174 515134 636618
rect 514514 600938 514546 601174
rect 514782 600938 514866 601174
rect 515102 600938 515134 601174
rect 514514 600854 515134 600938
rect 514514 600618 514546 600854
rect 514782 600618 514866 600854
rect 515102 600618 515134 600854
rect 514514 565174 515134 600618
rect 514514 564938 514546 565174
rect 514782 564938 514866 565174
rect 515102 564938 515134 565174
rect 514514 564854 515134 564938
rect 514514 564618 514546 564854
rect 514782 564618 514866 564854
rect 515102 564618 515134 564854
rect 514514 529174 515134 564618
rect 514514 528938 514546 529174
rect 514782 528938 514866 529174
rect 515102 528938 515134 529174
rect 514514 528854 515134 528938
rect 514514 528618 514546 528854
rect 514782 528618 514866 528854
rect 515102 528618 515134 528854
rect 514514 493174 515134 528618
rect 514514 492938 514546 493174
rect 514782 492938 514866 493174
rect 515102 492938 515134 493174
rect 514514 492854 515134 492938
rect 514514 492618 514546 492854
rect 514782 492618 514866 492854
rect 515102 492618 515134 492854
rect 514514 457174 515134 492618
rect 514514 456938 514546 457174
rect 514782 456938 514866 457174
rect 515102 456938 515134 457174
rect 514514 456854 515134 456938
rect 514514 456618 514546 456854
rect 514782 456618 514866 456854
rect 515102 456618 515134 456854
rect 514514 421174 515134 456618
rect 514514 420938 514546 421174
rect 514782 420938 514866 421174
rect 515102 420938 515134 421174
rect 514514 420854 515134 420938
rect 514514 420618 514546 420854
rect 514782 420618 514866 420854
rect 515102 420618 515134 420854
rect 514514 385174 515134 420618
rect 514514 384938 514546 385174
rect 514782 384938 514866 385174
rect 515102 384938 515134 385174
rect 514514 384854 515134 384938
rect 514514 384618 514546 384854
rect 514782 384618 514866 384854
rect 515102 384618 515134 384854
rect 514514 349174 515134 384618
rect 514514 348938 514546 349174
rect 514782 348938 514866 349174
rect 515102 348938 515134 349174
rect 514514 348854 515134 348938
rect 514514 348618 514546 348854
rect 514782 348618 514866 348854
rect 515102 348618 515134 348854
rect 514514 313174 515134 348618
rect 514514 312938 514546 313174
rect 514782 312938 514866 313174
rect 515102 312938 515134 313174
rect 514514 312854 515134 312938
rect 514514 312618 514546 312854
rect 514782 312618 514866 312854
rect 515102 312618 515134 312854
rect 514514 277174 515134 312618
rect 514514 276938 514546 277174
rect 514782 276938 514866 277174
rect 515102 276938 515134 277174
rect 514514 276854 515134 276938
rect 514514 276618 514546 276854
rect 514782 276618 514866 276854
rect 515102 276618 515134 276854
rect 514514 241174 515134 276618
rect 514514 240938 514546 241174
rect 514782 240938 514866 241174
rect 515102 240938 515134 241174
rect 514514 240854 515134 240938
rect 514514 240618 514546 240854
rect 514782 240618 514866 240854
rect 515102 240618 515134 240854
rect 514514 205174 515134 240618
rect 514514 204938 514546 205174
rect 514782 204938 514866 205174
rect 515102 204938 515134 205174
rect 514514 204854 515134 204938
rect 514514 204618 514546 204854
rect 514782 204618 514866 204854
rect 515102 204618 515134 204854
rect 514514 169174 515134 204618
rect 514514 168938 514546 169174
rect 514782 168938 514866 169174
rect 515102 168938 515134 169174
rect 514514 168854 515134 168938
rect 514514 168618 514546 168854
rect 514782 168618 514866 168854
rect 515102 168618 515134 168854
rect 514514 133174 515134 168618
rect 514514 132938 514546 133174
rect 514782 132938 514866 133174
rect 515102 132938 515134 133174
rect 514514 132854 515134 132938
rect 514514 132618 514546 132854
rect 514782 132618 514866 132854
rect 515102 132618 515134 132854
rect 514514 97174 515134 132618
rect 514514 96938 514546 97174
rect 514782 96938 514866 97174
rect 515102 96938 515134 97174
rect 514514 96854 515134 96938
rect 514514 96618 514546 96854
rect 514782 96618 514866 96854
rect 515102 96618 515134 96854
rect 514514 61174 515134 96618
rect 514514 60938 514546 61174
rect 514782 60938 514866 61174
rect 515102 60938 515134 61174
rect 514514 60854 515134 60938
rect 514514 60618 514546 60854
rect 514782 60618 514866 60854
rect 515102 60618 515134 60854
rect 514514 25174 515134 60618
rect 514514 24938 514546 25174
rect 514782 24938 514866 25174
rect 515102 24938 515134 25174
rect 514514 24854 515134 24938
rect 514514 24618 514546 24854
rect 514782 24618 514866 24854
rect 515102 24618 515134 24854
rect 514514 -3226 515134 24618
rect 514514 -3462 514546 -3226
rect 514782 -3462 514866 -3226
rect 515102 -3462 515134 -3226
rect 514514 -3546 515134 -3462
rect 514514 -3782 514546 -3546
rect 514782 -3782 514866 -3546
rect 515102 -3782 515134 -3546
rect 514514 -3814 515134 -3782
rect 518234 676894 518854 709082
rect 518234 676658 518266 676894
rect 518502 676658 518586 676894
rect 518822 676658 518854 676894
rect 518234 676574 518854 676658
rect 518234 676338 518266 676574
rect 518502 676338 518586 676574
rect 518822 676338 518854 676574
rect 518234 640894 518854 676338
rect 518234 640658 518266 640894
rect 518502 640658 518586 640894
rect 518822 640658 518854 640894
rect 518234 640574 518854 640658
rect 518234 640338 518266 640574
rect 518502 640338 518586 640574
rect 518822 640338 518854 640574
rect 518234 604894 518854 640338
rect 518234 604658 518266 604894
rect 518502 604658 518586 604894
rect 518822 604658 518854 604894
rect 518234 604574 518854 604658
rect 518234 604338 518266 604574
rect 518502 604338 518586 604574
rect 518822 604338 518854 604574
rect 518234 568894 518854 604338
rect 518234 568658 518266 568894
rect 518502 568658 518586 568894
rect 518822 568658 518854 568894
rect 518234 568574 518854 568658
rect 518234 568338 518266 568574
rect 518502 568338 518586 568574
rect 518822 568338 518854 568574
rect 518234 532894 518854 568338
rect 518234 532658 518266 532894
rect 518502 532658 518586 532894
rect 518822 532658 518854 532894
rect 518234 532574 518854 532658
rect 518234 532338 518266 532574
rect 518502 532338 518586 532574
rect 518822 532338 518854 532574
rect 518234 496894 518854 532338
rect 518234 496658 518266 496894
rect 518502 496658 518586 496894
rect 518822 496658 518854 496894
rect 518234 496574 518854 496658
rect 518234 496338 518266 496574
rect 518502 496338 518586 496574
rect 518822 496338 518854 496574
rect 518234 460894 518854 496338
rect 518234 460658 518266 460894
rect 518502 460658 518586 460894
rect 518822 460658 518854 460894
rect 518234 460574 518854 460658
rect 518234 460338 518266 460574
rect 518502 460338 518586 460574
rect 518822 460338 518854 460574
rect 518234 424894 518854 460338
rect 518234 424658 518266 424894
rect 518502 424658 518586 424894
rect 518822 424658 518854 424894
rect 518234 424574 518854 424658
rect 518234 424338 518266 424574
rect 518502 424338 518586 424574
rect 518822 424338 518854 424574
rect 518234 388894 518854 424338
rect 518234 388658 518266 388894
rect 518502 388658 518586 388894
rect 518822 388658 518854 388894
rect 518234 388574 518854 388658
rect 518234 388338 518266 388574
rect 518502 388338 518586 388574
rect 518822 388338 518854 388574
rect 518234 352894 518854 388338
rect 518234 352658 518266 352894
rect 518502 352658 518586 352894
rect 518822 352658 518854 352894
rect 518234 352574 518854 352658
rect 518234 352338 518266 352574
rect 518502 352338 518586 352574
rect 518822 352338 518854 352574
rect 518234 316894 518854 352338
rect 518234 316658 518266 316894
rect 518502 316658 518586 316894
rect 518822 316658 518854 316894
rect 518234 316574 518854 316658
rect 518234 316338 518266 316574
rect 518502 316338 518586 316574
rect 518822 316338 518854 316574
rect 518234 280894 518854 316338
rect 518234 280658 518266 280894
rect 518502 280658 518586 280894
rect 518822 280658 518854 280894
rect 518234 280574 518854 280658
rect 518234 280338 518266 280574
rect 518502 280338 518586 280574
rect 518822 280338 518854 280574
rect 518234 244894 518854 280338
rect 518234 244658 518266 244894
rect 518502 244658 518586 244894
rect 518822 244658 518854 244894
rect 518234 244574 518854 244658
rect 518234 244338 518266 244574
rect 518502 244338 518586 244574
rect 518822 244338 518854 244574
rect 518234 208894 518854 244338
rect 518234 208658 518266 208894
rect 518502 208658 518586 208894
rect 518822 208658 518854 208894
rect 518234 208574 518854 208658
rect 518234 208338 518266 208574
rect 518502 208338 518586 208574
rect 518822 208338 518854 208574
rect 518234 172894 518854 208338
rect 518234 172658 518266 172894
rect 518502 172658 518586 172894
rect 518822 172658 518854 172894
rect 518234 172574 518854 172658
rect 518234 172338 518266 172574
rect 518502 172338 518586 172574
rect 518822 172338 518854 172574
rect 518234 136894 518854 172338
rect 518234 136658 518266 136894
rect 518502 136658 518586 136894
rect 518822 136658 518854 136894
rect 518234 136574 518854 136658
rect 518234 136338 518266 136574
rect 518502 136338 518586 136574
rect 518822 136338 518854 136574
rect 518234 100894 518854 136338
rect 518234 100658 518266 100894
rect 518502 100658 518586 100894
rect 518822 100658 518854 100894
rect 518234 100574 518854 100658
rect 518234 100338 518266 100574
rect 518502 100338 518586 100574
rect 518822 100338 518854 100574
rect 518234 64894 518854 100338
rect 518234 64658 518266 64894
rect 518502 64658 518586 64894
rect 518822 64658 518854 64894
rect 518234 64574 518854 64658
rect 518234 64338 518266 64574
rect 518502 64338 518586 64574
rect 518822 64338 518854 64574
rect 518234 28894 518854 64338
rect 518234 28658 518266 28894
rect 518502 28658 518586 28894
rect 518822 28658 518854 28894
rect 518234 28574 518854 28658
rect 518234 28338 518266 28574
rect 518502 28338 518586 28574
rect 518822 28338 518854 28574
rect 518234 -5146 518854 28338
rect 520794 704838 521414 705830
rect 520794 704602 520826 704838
rect 521062 704602 521146 704838
rect 521382 704602 521414 704838
rect 520794 704518 521414 704602
rect 520794 704282 520826 704518
rect 521062 704282 521146 704518
rect 521382 704282 521414 704518
rect 520794 687454 521414 704282
rect 520794 687218 520826 687454
rect 521062 687218 521146 687454
rect 521382 687218 521414 687454
rect 520794 687134 521414 687218
rect 520794 686898 520826 687134
rect 521062 686898 521146 687134
rect 521382 686898 521414 687134
rect 520794 651454 521414 686898
rect 520794 651218 520826 651454
rect 521062 651218 521146 651454
rect 521382 651218 521414 651454
rect 520794 651134 521414 651218
rect 520794 650898 520826 651134
rect 521062 650898 521146 651134
rect 521382 650898 521414 651134
rect 520794 615454 521414 650898
rect 520794 615218 520826 615454
rect 521062 615218 521146 615454
rect 521382 615218 521414 615454
rect 520794 615134 521414 615218
rect 520794 614898 520826 615134
rect 521062 614898 521146 615134
rect 521382 614898 521414 615134
rect 520794 579454 521414 614898
rect 520794 579218 520826 579454
rect 521062 579218 521146 579454
rect 521382 579218 521414 579454
rect 520794 579134 521414 579218
rect 520794 578898 520826 579134
rect 521062 578898 521146 579134
rect 521382 578898 521414 579134
rect 520794 543454 521414 578898
rect 520794 543218 520826 543454
rect 521062 543218 521146 543454
rect 521382 543218 521414 543454
rect 520794 543134 521414 543218
rect 520794 542898 520826 543134
rect 521062 542898 521146 543134
rect 521382 542898 521414 543134
rect 520794 507454 521414 542898
rect 520794 507218 520826 507454
rect 521062 507218 521146 507454
rect 521382 507218 521414 507454
rect 520794 507134 521414 507218
rect 520794 506898 520826 507134
rect 521062 506898 521146 507134
rect 521382 506898 521414 507134
rect 520794 471454 521414 506898
rect 520794 471218 520826 471454
rect 521062 471218 521146 471454
rect 521382 471218 521414 471454
rect 520794 471134 521414 471218
rect 520794 470898 520826 471134
rect 521062 470898 521146 471134
rect 521382 470898 521414 471134
rect 520794 435454 521414 470898
rect 520794 435218 520826 435454
rect 521062 435218 521146 435454
rect 521382 435218 521414 435454
rect 520794 435134 521414 435218
rect 520794 434898 520826 435134
rect 521062 434898 521146 435134
rect 521382 434898 521414 435134
rect 520794 399454 521414 434898
rect 520794 399218 520826 399454
rect 521062 399218 521146 399454
rect 521382 399218 521414 399454
rect 520794 399134 521414 399218
rect 520794 398898 520826 399134
rect 521062 398898 521146 399134
rect 521382 398898 521414 399134
rect 520794 363454 521414 398898
rect 520794 363218 520826 363454
rect 521062 363218 521146 363454
rect 521382 363218 521414 363454
rect 520794 363134 521414 363218
rect 520794 362898 520826 363134
rect 521062 362898 521146 363134
rect 521382 362898 521414 363134
rect 520794 327454 521414 362898
rect 520794 327218 520826 327454
rect 521062 327218 521146 327454
rect 521382 327218 521414 327454
rect 520794 327134 521414 327218
rect 520794 326898 520826 327134
rect 521062 326898 521146 327134
rect 521382 326898 521414 327134
rect 520794 291454 521414 326898
rect 520794 291218 520826 291454
rect 521062 291218 521146 291454
rect 521382 291218 521414 291454
rect 520794 291134 521414 291218
rect 520794 290898 520826 291134
rect 521062 290898 521146 291134
rect 521382 290898 521414 291134
rect 520794 255454 521414 290898
rect 520794 255218 520826 255454
rect 521062 255218 521146 255454
rect 521382 255218 521414 255454
rect 520794 255134 521414 255218
rect 520794 254898 520826 255134
rect 521062 254898 521146 255134
rect 521382 254898 521414 255134
rect 520794 219454 521414 254898
rect 520794 219218 520826 219454
rect 521062 219218 521146 219454
rect 521382 219218 521414 219454
rect 520794 219134 521414 219218
rect 520794 218898 520826 219134
rect 521062 218898 521146 219134
rect 521382 218898 521414 219134
rect 520794 183454 521414 218898
rect 520794 183218 520826 183454
rect 521062 183218 521146 183454
rect 521382 183218 521414 183454
rect 520794 183134 521414 183218
rect 520794 182898 520826 183134
rect 521062 182898 521146 183134
rect 521382 182898 521414 183134
rect 520794 147454 521414 182898
rect 520794 147218 520826 147454
rect 521062 147218 521146 147454
rect 521382 147218 521414 147454
rect 520794 147134 521414 147218
rect 520794 146898 520826 147134
rect 521062 146898 521146 147134
rect 521382 146898 521414 147134
rect 520794 111454 521414 146898
rect 520794 111218 520826 111454
rect 521062 111218 521146 111454
rect 521382 111218 521414 111454
rect 520794 111134 521414 111218
rect 520794 110898 520826 111134
rect 521062 110898 521146 111134
rect 521382 110898 521414 111134
rect 520794 75454 521414 110898
rect 520794 75218 520826 75454
rect 521062 75218 521146 75454
rect 521382 75218 521414 75454
rect 520794 75134 521414 75218
rect 520794 74898 520826 75134
rect 521062 74898 521146 75134
rect 521382 74898 521414 75134
rect 520794 39454 521414 74898
rect 520794 39218 520826 39454
rect 521062 39218 521146 39454
rect 521382 39218 521414 39454
rect 520794 39134 521414 39218
rect 520794 38898 520826 39134
rect 521062 38898 521146 39134
rect 521382 38898 521414 39134
rect 520794 3454 521414 38898
rect 520794 3218 520826 3454
rect 521062 3218 521146 3454
rect 521382 3218 521414 3454
rect 520794 3134 521414 3218
rect 520794 2898 520826 3134
rect 521062 2898 521146 3134
rect 521382 2898 521414 3134
rect 520794 -346 521414 2898
rect 520794 -582 520826 -346
rect 521062 -582 521146 -346
rect 521382 -582 521414 -346
rect 520794 -666 521414 -582
rect 520794 -902 520826 -666
rect 521062 -902 521146 -666
rect 521382 -902 521414 -666
rect 520794 -1894 521414 -902
rect 521954 680614 522574 711002
rect 531954 710598 532574 711590
rect 531954 710362 531986 710598
rect 532222 710362 532306 710598
rect 532542 710362 532574 710598
rect 531954 710278 532574 710362
rect 531954 710042 531986 710278
rect 532222 710042 532306 710278
rect 532542 710042 532574 710278
rect 528234 708678 528854 709670
rect 528234 708442 528266 708678
rect 528502 708442 528586 708678
rect 528822 708442 528854 708678
rect 528234 708358 528854 708442
rect 528234 708122 528266 708358
rect 528502 708122 528586 708358
rect 528822 708122 528854 708358
rect 521954 680378 521986 680614
rect 522222 680378 522306 680614
rect 522542 680378 522574 680614
rect 521954 680294 522574 680378
rect 521954 680058 521986 680294
rect 522222 680058 522306 680294
rect 522542 680058 522574 680294
rect 521954 644614 522574 680058
rect 521954 644378 521986 644614
rect 522222 644378 522306 644614
rect 522542 644378 522574 644614
rect 521954 644294 522574 644378
rect 521954 644058 521986 644294
rect 522222 644058 522306 644294
rect 522542 644058 522574 644294
rect 521954 608614 522574 644058
rect 521954 608378 521986 608614
rect 522222 608378 522306 608614
rect 522542 608378 522574 608614
rect 521954 608294 522574 608378
rect 521954 608058 521986 608294
rect 522222 608058 522306 608294
rect 522542 608058 522574 608294
rect 521954 572614 522574 608058
rect 521954 572378 521986 572614
rect 522222 572378 522306 572614
rect 522542 572378 522574 572614
rect 521954 572294 522574 572378
rect 521954 572058 521986 572294
rect 522222 572058 522306 572294
rect 522542 572058 522574 572294
rect 521954 536614 522574 572058
rect 521954 536378 521986 536614
rect 522222 536378 522306 536614
rect 522542 536378 522574 536614
rect 521954 536294 522574 536378
rect 521954 536058 521986 536294
rect 522222 536058 522306 536294
rect 522542 536058 522574 536294
rect 521954 500614 522574 536058
rect 521954 500378 521986 500614
rect 522222 500378 522306 500614
rect 522542 500378 522574 500614
rect 521954 500294 522574 500378
rect 521954 500058 521986 500294
rect 522222 500058 522306 500294
rect 522542 500058 522574 500294
rect 521954 464614 522574 500058
rect 521954 464378 521986 464614
rect 522222 464378 522306 464614
rect 522542 464378 522574 464614
rect 521954 464294 522574 464378
rect 521954 464058 521986 464294
rect 522222 464058 522306 464294
rect 522542 464058 522574 464294
rect 521954 428614 522574 464058
rect 521954 428378 521986 428614
rect 522222 428378 522306 428614
rect 522542 428378 522574 428614
rect 521954 428294 522574 428378
rect 521954 428058 521986 428294
rect 522222 428058 522306 428294
rect 522542 428058 522574 428294
rect 521954 392614 522574 428058
rect 521954 392378 521986 392614
rect 522222 392378 522306 392614
rect 522542 392378 522574 392614
rect 521954 392294 522574 392378
rect 521954 392058 521986 392294
rect 522222 392058 522306 392294
rect 522542 392058 522574 392294
rect 521954 356614 522574 392058
rect 521954 356378 521986 356614
rect 522222 356378 522306 356614
rect 522542 356378 522574 356614
rect 521954 356294 522574 356378
rect 521954 356058 521986 356294
rect 522222 356058 522306 356294
rect 522542 356058 522574 356294
rect 521954 320614 522574 356058
rect 521954 320378 521986 320614
rect 522222 320378 522306 320614
rect 522542 320378 522574 320614
rect 521954 320294 522574 320378
rect 521954 320058 521986 320294
rect 522222 320058 522306 320294
rect 522542 320058 522574 320294
rect 521954 284614 522574 320058
rect 521954 284378 521986 284614
rect 522222 284378 522306 284614
rect 522542 284378 522574 284614
rect 521954 284294 522574 284378
rect 521954 284058 521986 284294
rect 522222 284058 522306 284294
rect 522542 284058 522574 284294
rect 521954 248614 522574 284058
rect 521954 248378 521986 248614
rect 522222 248378 522306 248614
rect 522542 248378 522574 248614
rect 521954 248294 522574 248378
rect 521954 248058 521986 248294
rect 522222 248058 522306 248294
rect 522542 248058 522574 248294
rect 521954 212614 522574 248058
rect 521954 212378 521986 212614
rect 522222 212378 522306 212614
rect 522542 212378 522574 212614
rect 521954 212294 522574 212378
rect 521954 212058 521986 212294
rect 522222 212058 522306 212294
rect 522542 212058 522574 212294
rect 521954 176614 522574 212058
rect 521954 176378 521986 176614
rect 522222 176378 522306 176614
rect 522542 176378 522574 176614
rect 521954 176294 522574 176378
rect 521954 176058 521986 176294
rect 522222 176058 522306 176294
rect 522542 176058 522574 176294
rect 521954 140614 522574 176058
rect 521954 140378 521986 140614
rect 522222 140378 522306 140614
rect 522542 140378 522574 140614
rect 521954 140294 522574 140378
rect 521954 140058 521986 140294
rect 522222 140058 522306 140294
rect 522542 140058 522574 140294
rect 521954 104614 522574 140058
rect 521954 104378 521986 104614
rect 522222 104378 522306 104614
rect 522542 104378 522574 104614
rect 521954 104294 522574 104378
rect 521954 104058 521986 104294
rect 522222 104058 522306 104294
rect 522542 104058 522574 104294
rect 521954 68614 522574 104058
rect 521954 68378 521986 68614
rect 522222 68378 522306 68614
rect 522542 68378 522574 68614
rect 521954 68294 522574 68378
rect 521954 68058 521986 68294
rect 522222 68058 522306 68294
rect 522542 68058 522574 68294
rect 521954 32614 522574 68058
rect 521954 32378 521986 32614
rect 522222 32378 522306 32614
rect 522542 32378 522574 32614
rect 521954 32294 522574 32378
rect 521954 32058 521986 32294
rect 522222 32058 522306 32294
rect 522542 32058 522574 32294
rect 518234 -5382 518266 -5146
rect 518502 -5382 518586 -5146
rect 518822 -5382 518854 -5146
rect 518234 -5466 518854 -5382
rect 518234 -5702 518266 -5466
rect 518502 -5702 518586 -5466
rect 518822 -5702 518854 -5466
rect 518234 -5734 518854 -5702
rect 511954 -6342 511986 -6106
rect 512222 -6342 512306 -6106
rect 512542 -6342 512574 -6106
rect 511954 -6426 512574 -6342
rect 511954 -6662 511986 -6426
rect 512222 -6662 512306 -6426
rect 512542 -6662 512574 -6426
rect 511954 -7654 512574 -6662
rect 521954 -7066 522574 32058
rect 524514 706758 525134 707750
rect 524514 706522 524546 706758
rect 524782 706522 524866 706758
rect 525102 706522 525134 706758
rect 524514 706438 525134 706522
rect 524514 706202 524546 706438
rect 524782 706202 524866 706438
rect 525102 706202 525134 706438
rect 524514 691174 525134 706202
rect 524514 690938 524546 691174
rect 524782 690938 524866 691174
rect 525102 690938 525134 691174
rect 524514 690854 525134 690938
rect 524514 690618 524546 690854
rect 524782 690618 524866 690854
rect 525102 690618 525134 690854
rect 524514 655174 525134 690618
rect 524514 654938 524546 655174
rect 524782 654938 524866 655174
rect 525102 654938 525134 655174
rect 524514 654854 525134 654938
rect 524514 654618 524546 654854
rect 524782 654618 524866 654854
rect 525102 654618 525134 654854
rect 524514 619174 525134 654618
rect 524514 618938 524546 619174
rect 524782 618938 524866 619174
rect 525102 618938 525134 619174
rect 524514 618854 525134 618938
rect 524514 618618 524546 618854
rect 524782 618618 524866 618854
rect 525102 618618 525134 618854
rect 524514 583174 525134 618618
rect 524514 582938 524546 583174
rect 524782 582938 524866 583174
rect 525102 582938 525134 583174
rect 524514 582854 525134 582938
rect 524514 582618 524546 582854
rect 524782 582618 524866 582854
rect 525102 582618 525134 582854
rect 524514 547174 525134 582618
rect 524514 546938 524546 547174
rect 524782 546938 524866 547174
rect 525102 546938 525134 547174
rect 524514 546854 525134 546938
rect 524514 546618 524546 546854
rect 524782 546618 524866 546854
rect 525102 546618 525134 546854
rect 524514 511174 525134 546618
rect 524514 510938 524546 511174
rect 524782 510938 524866 511174
rect 525102 510938 525134 511174
rect 524514 510854 525134 510938
rect 524514 510618 524546 510854
rect 524782 510618 524866 510854
rect 525102 510618 525134 510854
rect 524514 475174 525134 510618
rect 524514 474938 524546 475174
rect 524782 474938 524866 475174
rect 525102 474938 525134 475174
rect 524514 474854 525134 474938
rect 524514 474618 524546 474854
rect 524782 474618 524866 474854
rect 525102 474618 525134 474854
rect 524514 439174 525134 474618
rect 524514 438938 524546 439174
rect 524782 438938 524866 439174
rect 525102 438938 525134 439174
rect 524514 438854 525134 438938
rect 524514 438618 524546 438854
rect 524782 438618 524866 438854
rect 525102 438618 525134 438854
rect 524514 403174 525134 438618
rect 524514 402938 524546 403174
rect 524782 402938 524866 403174
rect 525102 402938 525134 403174
rect 524514 402854 525134 402938
rect 524514 402618 524546 402854
rect 524782 402618 524866 402854
rect 525102 402618 525134 402854
rect 524514 367174 525134 402618
rect 524514 366938 524546 367174
rect 524782 366938 524866 367174
rect 525102 366938 525134 367174
rect 524514 366854 525134 366938
rect 524514 366618 524546 366854
rect 524782 366618 524866 366854
rect 525102 366618 525134 366854
rect 524514 331174 525134 366618
rect 524514 330938 524546 331174
rect 524782 330938 524866 331174
rect 525102 330938 525134 331174
rect 524514 330854 525134 330938
rect 524514 330618 524546 330854
rect 524782 330618 524866 330854
rect 525102 330618 525134 330854
rect 524514 295174 525134 330618
rect 524514 294938 524546 295174
rect 524782 294938 524866 295174
rect 525102 294938 525134 295174
rect 524514 294854 525134 294938
rect 524514 294618 524546 294854
rect 524782 294618 524866 294854
rect 525102 294618 525134 294854
rect 524514 259174 525134 294618
rect 524514 258938 524546 259174
rect 524782 258938 524866 259174
rect 525102 258938 525134 259174
rect 524514 258854 525134 258938
rect 524514 258618 524546 258854
rect 524782 258618 524866 258854
rect 525102 258618 525134 258854
rect 524514 223174 525134 258618
rect 524514 222938 524546 223174
rect 524782 222938 524866 223174
rect 525102 222938 525134 223174
rect 524514 222854 525134 222938
rect 524514 222618 524546 222854
rect 524782 222618 524866 222854
rect 525102 222618 525134 222854
rect 524514 187174 525134 222618
rect 524514 186938 524546 187174
rect 524782 186938 524866 187174
rect 525102 186938 525134 187174
rect 524514 186854 525134 186938
rect 524514 186618 524546 186854
rect 524782 186618 524866 186854
rect 525102 186618 525134 186854
rect 524514 151174 525134 186618
rect 524514 150938 524546 151174
rect 524782 150938 524866 151174
rect 525102 150938 525134 151174
rect 524514 150854 525134 150938
rect 524514 150618 524546 150854
rect 524782 150618 524866 150854
rect 525102 150618 525134 150854
rect 524514 115174 525134 150618
rect 524514 114938 524546 115174
rect 524782 114938 524866 115174
rect 525102 114938 525134 115174
rect 524514 114854 525134 114938
rect 524514 114618 524546 114854
rect 524782 114618 524866 114854
rect 525102 114618 525134 114854
rect 524514 79174 525134 114618
rect 524514 78938 524546 79174
rect 524782 78938 524866 79174
rect 525102 78938 525134 79174
rect 524514 78854 525134 78938
rect 524514 78618 524546 78854
rect 524782 78618 524866 78854
rect 525102 78618 525134 78854
rect 524514 43174 525134 78618
rect 524514 42938 524546 43174
rect 524782 42938 524866 43174
rect 525102 42938 525134 43174
rect 524514 42854 525134 42938
rect 524514 42618 524546 42854
rect 524782 42618 524866 42854
rect 525102 42618 525134 42854
rect 524514 7174 525134 42618
rect 524514 6938 524546 7174
rect 524782 6938 524866 7174
rect 525102 6938 525134 7174
rect 524514 6854 525134 6938
rect 524514 6618 524546 6854
rect 524782 6618 524866 6854
rect 525102 6618 525134 6854
rect 524514 -2266 525134 6618
rect 524514 -2502 524546 -2266
rect 524782 -2502 524866 -2266
rect 525102 -2502 525134 -2266
rect 524514 -2586 525134 -2502
rect 524514 -2822 524546 -2586
rect 524782 -2822 524866 -2586
rect 525102 -2822 525134 -2586
rect 524514 -3814 525134 -2822
rect 528234 694894 528854 708122
rect 528234 694658 528266 694894
rect 528502 694658 528586 694894
rect 528822 694658 528854 694894
rect 528234 694574 528854 694658
rect 528234 694338 528266 694574
rect 528502 694338 528586 694574
rect 528822 694338 528854 694574
rect 528234 658894 528854 694338
rect 528234 658658 528266 658894
rect 528502 658658 528586 658894
rect 528822 658658 528854 658894
rect 528234 658574 528854 658658
rect 528234 658338 528266 658574
rect 528502 658338 528586 658574
rect 528822 658338 528854 658574
rect 528234 622894 528854 658338
rect 528234 622658 528266 622894
rect 528502 622658 528586 622894
rect 528822 622658 528854 622894
rect 528234 622574 528854 622658
rect 528234 622338 528266 622574
rect 528502 622338 528586 622574
rect 528822 622338 528854 622574
rect 528234 586894 528854 622338
rect 528234 586658 528266 586894
rect 528502 586658 528586 586894
rect 528822 586658 528854 586894
rect 528234 586574 528854 586658
rect 528234 586338 528266 586574
rect 528502 586338 528586 586574
rect 528822 586338 528854 586574
rect 528234 550894 528854 586338
rect 528234 550658 528266 550894
rect 528502 550658 528586 550894
rect 528822 550658 528854 550894
rect 528234 550574 528854 550658
rect 528234 550338 528266 550574
rect 528502 550338 528586 550574
rect 528822 550338 528854 550574
rect 528234 514894 528854 550338
rect 528234 514658 528266 514894
rect 528502 514658 528586 514894
rect 528822 514658 528854 514894
rect 528234 514574 528854 514658
rect 528234 514338 528266 514574
rect 528502 514338 528586 514574
rect 528822 514338 528854 514574
rect 528234 478894 528854 514338
rect 528234 478658 528266 478894
rect 528502 478658 528586 478894
rect 528822 478658 528854 478894
rect 528234 478574 528854 478658
rect 528234 478338 528266 478574
rect 528502 478338 528586 478574
rect 528822 478338 528854 478574
rect 528234 442894 528854 478338
rect 528234 442658 528266 442894
rect 528502 442658 528586 442894
rect 528822 442658 528854 442894
rect 528234 442574 528854 442658
rect 528234 442338 528266 442574
rect 528502 442338 528586 442574
rect 528822 442338 528854 442574
rect 528234 406894 528854 442338
rect 528234 406658 528266 406894
rect 528502 406658 528586 406894
rect 528822 406658 528854 406894
rect 528234 406574 528854 406658
rect 528234 406338 528266 406574
rect 528502 406338 528586 406574
rect 528822 406338 528854 406574
rect 528234 370894 528854 406338
rect 528234 370658 528266 370894
rect 528502 370658 528586 370894
rect 528822 370658 528854 370894
rect 528234 370574 528854 370658
rect 528234 370338 528266 370574
rect 528502 370338 528586 370574
rect 528822 370338 528854 370574
rect 528234 334894 528854 370338
rect 528234 334658 528266 334894
rect 528502 334658 528586 334894
rect 528822 334658 528854 334894
rect 528234 334574 528854 334658
rect 528234 334338 528266 334574
rect 528502 334338 528586 334574
rect 528822 334338 528854 334574
rect 528234 298894 528854 334338
rect 528234 298658 528266 298894
rect 528502 298658 528586 298894
rect 528822 298658 528854 298894
rect 528234 298574 528854 298658
rect 528234 298338 528266 298574
rect 528502 298338 528586 298574
rect 528822 298338 528854 298574
rect 528234 262894 528854 298338
rect 528234 262658 528266 262894
rect 528502 262658 528586 262894
rect 528822 262658 528854 262894
rect 528234 262574 528854 262658
rect 528234 262338 528266 262574
rect 528502 262338 528586 262574
rect 528822 262338 528854 262574
rect 528234 226894 528854 262338
rect 528234 226658 528266 226894
rect 528502 226658 528586 226894
rect 528822 226658 528854 226894
rect 528234 226574 528854 226658
rect 528234 226338 528266 226574
rect 528502 226338 528586 226574
rect 528822 226338 528854 226574
rect 528234 190894 528854 226338
rect 528234 190658 528266 190894
rect 528502 190658 528586 190894
rect 528822 190658 528854 190894
rect 528234 190574 528854 190658
rect 528234 190338 528266 190574
rect 528502 190338 528586 190574
rect 528822 190338 528854 190574
rect 528234 154894 528854 190338
rect 528234 154658 528266 154894
rect 528502 154658 528586 154894
rect 528822 154658 528854 154894
rect 528234 154574 528854 154658
rect 528234 154338 528266 154574
rect 528502 154338 528586 154574
rect 528822 154338 528854 154574
rect 528234 118894 528854 154338
rect 528234 118658 528266 118894
rect 528502 118658 528586 118894
rect 528822 118658 528854 118894
rect 528234 118574 528854 118658
rect 528234 118338 528266 118574
rect 528502 118338 528586 118574
rect 528822 118338 528854 118574
rect 528234 82894 528854 118338
rect 528234 82658 528266 82894
rect 528502 82658 528586 82894
rect 528822 82658 528854 82894
rect 528234 82574 528854 82658
rect 528234 82338 528266 82574
rect 528502 82338 528586 82574
rect 528822 82338 528854 82574
rect 528234 46894 528854 82338
rect 528234 46658 528266 46894
rect 528502 46658 528586 46894
rect 528822 46658 528854 46894
rect 528234 46574 528854 46658
rect 528234 46338 528266 46574
rect 528502 46338 528586 46574
rect 528822 46338 528854 46574
rect 528234 10894 528854 46338
rect 528234 10658 528266 10894
rect 528502 10658 528586 10894
rect 528822 10658 528854 10894
rect 528234 10574 528854 10658
rect 528234 10338 528266 10574
rect 528502 10338 528586 10574
rect 528822 10338 528854 10574
rect 528234 -4186 528854 10338
rect 530794 705798 531414 705830
rect 530794 705562 530826 705798
rect 531062 705562 531146 705798
rect 531382 705562 531414 705798
rect 530794 705478 531414 705562
rect 530794 705242 530826 705478
rect 531062 705242 531146 705478
rect 531382 705242 531414 705478
rect 530794 669454 531414 705242
rect 530794 669218 530826 669454
rect 531062 669218 531146 669454
rect 531382 669218 531414 669454
rect 530794 669134 531414 669218
rect 530794 668898 530826 669134
rect 531062 668898 531146 669134
rect 531382 668898 531414 669134
rect 530794 633454 531414 668898
rect 530794 633218 530826 633454
rect 531062 633218 531146 633454
rect 531382 633218 531414 633454
rect 530794 633134 531414 633218
rect 530794 632898 530826 633134
rect 531062 632898 531146 633134
rect 531382 632898 531414 633134
rect 530794 597454 531414 632898
rect 530794 597218 530826 597454
rect 531062 597218 531146 597454
rect 531382 597218 531414 597454
rect 530794 597134 531414 597218
rect 530794 596898 530826 597134
rect 531062 596898 531146 597134
rect 531382 596898 531414 597134
rect 530794 561454 531414 596898
rect 530794 561218 530826 561454
rect 531062 561218 531146 561454
rect 531382 561218 531414 561454
rect 530794 561134 531414 561218
rect 530794 560898 530826 561134
rect 531062 560898 531146 561134
rect 531382 560898 531414 561134
rect 530794 525454 531414 560898
rect 530794 525218 530826 525454
rect 531062 525218 531146 525454
rect 531382 525218 531414 525454
rect 530794 525134 531414 525218
rect 530794 524898 530826 525134
rect 531062 524898 531146 525134
rect 531382 524898 531414 525134
rect 530794 489454 531414 524898
rect 530794 489218 530826 489454
rect 531062 489218 531146 489454
rect 531382 489218 531414 489454
rect 530794 489134 531414 489218
rect 530794 488898 530826 489134
rect 531062 488898 531146 489134
rect 531382 488898 531414 489134
rect 530794 453454 531414 488898
rect 530794 453218 530826 453454
rect 531062 453218 531146 453454
rect 531382 453218 531414 453454
rect 530794 453134 531414 453218
rect 530794 452898 530826 453134
rect 531062 452898 531146 453134
rect 531382 452898 531414 453134
rect 530794 417454 531414 452898
rect 530794 417218 530826 417454
rect 531062 417218 531146 417454
rect 531382 417218 531414 417454
rect 530794 417134 531414 417218
rect 530794 416898 530826 417134
rect 531062 416898 531146 417134
rect 531382 416898 531414 417134
rect 530794 381454 531414 416898
rect 530794 381218 530826 381454
rect 531062 381218 531146 381454
rect 531382 381218 531414 381454
rect 530794 381134 531414 381218
rect 530794 380898 530826 381134
rect 531062 380898 531146 381134
rect 531382 380898 531414 381134
rect 530794 345454 531414 380898
rect 530794 345218 530826 345454
rect 531062 345218 531146 345454
rect 531382 345218 531414 345454
rect 530794 345134 531414 345218
rect 530794 344898 530826 345134
rect 531062 344898 531146 345134
rect 531382 344898 531414 345134
rect 530794 309454 531414 344898
rect 530794 309218 530826 309454
rect 531062 309218 531146 309454
rect 531382 309218 531414 309454
rect 530794 309134 531414 309218
rect 530794 308898 530826 309134
rect 531062 308898 531146 309134
rect 531382 308898 531414 309134
rect 530794 273454 531414 308898
rect 530794 273218 530826 273454
rect 531062 273218 531146 273454
rect 531382 273218 531414 273454
rect 530794 273134 531414 273218
rect 530794 272898 530826 273134
rect 531062 272898 531146 273134
rect 531382 272898 531414 273134
rect 530794 237454 531414 272898
rect 530794 237218 530826 237454
rect 531062 237218 531146 237454
rect 531382 237218 531414 237454
rect 530794 237134 531414 237218
rect 530794 236898 530826 237134
rect 531062 236898 531146 237134
rect 531382 236898 531414 237134
rect 530794 201454 531414 236898
rect 530794 201218 530826 201454
rect 531062 201218 531146 201454
rect 531382 201218 531414 201454
rect 530794 201134 531414 201218
rect 530794 200898 530826 201134
rect 531062 200898 531146 201134
rect 531382 200898 531414 201134
rect 530794 165454 531414 200898
rect 530794 165218 530826 165454
rect 531062 165218 531146 165454
rect 531382 165218 531414 165454
rect 530794 165134 531414 165218
rect 530794 164898 530826 165134
rect 531062 164898 531146 165134
rect 531382 164898 531414 165134
rect 530794 129454 531414 164898
rect 530794 129218 530826 129454
rect 531062 129218 531146 129454
rect 531382 129218 531414 129454
rect 530794 129134 531414 129218
rect 530794 128898 530826 129134
rect 531062 128898 531146 129134
rect 531382 128898 531414 129134
rect 530794 93454 531414 128898
rect 530794 93218 530826 93454
rect 531062 93218 531146 93454
rect 531382 93218 531414 93454
rect 530794 93134 531414 93218
rect 530794 92898 530826 93134
rect 531062 92898 531146 93134
rect 531382 92898 531414 93134
rect 530794 57454 531414 92898
rect 530794 57218 530826 57454
rect 531062 57218 531146 57454
rect 531382 57218 531414 57454
rect 530794 57134 531414 57218
rect 530794 56898 530826 57134
rect 531062 56898 531146 57134
rect 531382 56898 531414 57134
rect 530794 21454 531414 56898
rect 530794 21218 530826 21454
rect 531062 21218 531146 21454
rect 531382 21218 531414 21454
rect 530794 21134 531414 21218
rect 530794 20898 530826 21134
rect 531062 20898 531146 21134
rect 531382 20898 531414 21134
rect 530794 -1306 531414 20898
rect 530794 -1542 530826 -1306
rect 531062 -1542 531146 -1306
rect 531382 -1542 531414 -1306
rect 530794 -1626 531414 -1542
rect 530794 -1862 530826 -1626
rect 531062 -1862 531146 -1626
rect 531382 -1862 531414 -1626
rect 530794 -1894 531414 -1862
rect 531954 698614 532574 710042
rect 541954 711558 542574 711590
rect 541954 711322 541986 711558
rect 542222 711322 542306 711558
rect 542542 711322 542574 711558
rect 541954 711238 542574 711322
rect 541954 711002 541986 711238
rect 542222 711002 542306 711238
rect 542542 711002 542574 711238
rect 538234 709638 538854 709670
rect 538234 709402 538266 709638
rect 538502 709402 538586 709638
rect 538822 709402 538854 709638
rect 538234 709318 538854 709402
rect 538234 709082 538266 709318
rect 538502 709082 538586 709318
rect 538822 709082 538854 709318
rect 531954 698378 531986 698614
rect 532222 698378 532306 698614
rect 532542 698378 532574 698614
rect 531954 698294 532574 698378
rect 531954 698058 531986 698294
rect 532222 698058 532306 698294
rect 532542 698058 532574 698294
rect 531954 662614 532574 698058
rect 531954 662378 531986 662614
rect 532222 662378 532306 662614
rect 532542 662378 532574 662614
rect 531954 662294 532574 662378
rect 531954 662058 531986 662294
rect 532222 662058 532306 662294
rect 532542 662058 532574 662294
rect 531954 626614 532574 662058
rect 531954 626378 531986 626614
rect 532222 626378 532306 626614
rect 532542 626378 532574 626614
rect 531954 626294 532574 626378
rect 531954 626058 531986 626294
rect 532222 626058 532306 626294
rect 532542 626058 532574 626294
rect 531954 590614 532574 626058
rect 531954 590378 531986 590614
rect 532222 590378 532306 590614
rect 532542 590378 532574 590614
rect 531954 590294 532574 590378
rect 531954 590058 531986 590294
rect 532222 590058 532306 590294
rect 532542 590058 532574 590294
rect 531954 554614 532574 590058
rect 531954 554378 531986 554614
rect 532222 554378 532306 554614
rect 532542 554378 532574 554614
rect 531954 554294 532574 554378
rect 531954 554058 531986 554294
rect 532222 554058 532306 554294
rect 532542 554058 532574 554294
rect 531954 518614 532574 554058
rect 531954 518378 531986 518614
rect 532222 518378 532306 518614
rect 532542 518378 532574 518614
rect 531954 518294 532574 518378
rect 531954 518058 531986 518294
rect 532222 518058 532306 518294
rect 532542 518058 532574 518294
rect 531954 482614 532574 518058
rect 531954 482378 531986 482614
rect 532222 482378 532306 482614
rect 532542 482378 532574 482614
rect 531954 482294 532574 482378
rect 531954 482058 531986 482294
rect 532222 482058 532306 482294
rect 532542 482058 532574 482294
rect 531954 446614 532574 482058
rect 531954 446378 531986 446614
rect 532222 446378 532306 446614
rect 532542 446378 532574 446614
rect 531954 446294 532574 446378
rect 531954 446058 531986 446294
rect 532222 446058 532306 446294
rect 532542 446058 532574 446294
rect 531954 410614 532574 446058
rect 531954 410378 531986 410614
rect 532222 410378 532306 410614
rect 532542 410378 532574 410614
rect 531954 410294 532574 410378
rect 531954 410058 531986 410294
rect 532222 410058 532306 410294
rect 532542 410058 532574 410294
rect 531954 374614 532574 410058
rect 531954 374378 531986 374614
rect 532222 374378 532306 374614
rect 532542 374378 532574 374614
rect 531954 374294 532574 374378
rect 531954 374058 531986 374294
rect 532222 374058 532306 374294
rect 532542 374058 532574 374294
rect 531954 338614 532574 374058
rect 531954 338378 531986 338614
rect 532222 338378 532306 338614
rect 532542 338378 532574 338614
rect 531954 338294 532574 338378
rect 531954 338058 531986 338294
rect 532222 338058 532306 338294
rect 532542 338058 532574 338294
rect 531954 302614 532574 338058
rect 531954 302378 531986 302614
rect 532222 302378 532306 302614
rect 532542 302378 532574 302614
rect 531954 302294 532574 302378
rect 531954 302058 531986 302294
rect 532222 302058 532306 302294
rect 532542 302058 532574 302294
rect 531954 266614 532574 302058
rect 531954 266378 531986 266614
rect 532222 266378 532306 266614
rect 532542 266378 532574 266614
rect 531954 266294 532574 266378
rect 531954 266058 531986 266294
rect 532222 266058 532306 266294
rect 532542 266058 532574 266294
rect 531954 230614 532574 266058
rect 531954 230378 531986 230614
rect 532222 230378 532306 230614
rect 532542 230378 532574 230614
rect 531954 230294 532574 230378
rect 531954 230058 531986 230294
rect 532222 230058 532306 230294
rect 532542 230058 532574 230294
rect 531954 194614 532574 230058
rect 531954 194378 531986 194614
rect 532222 194378 532306 194614
rect 532542 194378 532574 194614
rect 531954 194294 532574 194378
rect 531954 194058 531986 194294
rect 532222 194058 532306 194294
rect 532542 194058 532574 194294
rect 531954 158614 532574 194058
rect 531954 158378 531986 158614
rect 532222 158378 532306 158614
rect 532542 158378 532574 158614
rect 531954 158294 532574 158378
rect 531954 158058 531986 158294
rect 532222 158058 532306 158294
rect 532542 158058 532574 158294
rect 531954 122614 532574 158058
rect 531954 122378 531986 122614
rect 532222 122378 532306 122614
rect 532542 122378 532574 122614
rect 531954 122294 532574 122378
rect 531954 122058 531986 122294
rect 532222 122058 532306 122294
rect 532542 122058 532574 122294
rect 531954 86614 532574 122058
rect 531954 86378 531986 86614
rect 532222 86378 532306 86614
rect 532542 86378 532574 86614
rect 531954 86294 532574 86378
rect 531954 86058 531986 86294
rect 532222 86058 532306 86294
rect 532542 86058 532574 86294
rect 531954 50614 532574 86058
rect 531954 50378 531986 50614
rect 532222 50378 532306 50614
rect 532542 50378 532574 50614
rect 531954 50294 532574 50378
rect 531954 50058 531986 50294
rect 532222 50058 532306 50294
rect 532542 50058 532574 50294
rect 531954 14614 532574 50058
rect 531954 14378 531986 14614
rect 532222 14378 532306 14614
rect 532542 14378 532574 14614
rect 531954 14294 532574 14378
rect 531954 14058 531986 14294
rect 532222 14058 532306 14294
rect 532542 14058 532574 14294
rect 528234 -4422 528266 -4186
rect 528502 -4422 528586 -4186
rect 528822 -4422 528854 -4186
rect 528234 -4506 528854 -4422
rect 528234 -4742 528266 -4506
rect 528502 -4742 528586 -4506
rect 528822 -4742 528854 -4506
rect 528234 -5734 528854 -4742
rect 521954 -7302 521986 -7066
rect 522222 -7302 522306 -7066
rect 522542 -7302 522574 -7066
rect 521954 -7386 522574 -7302
rect 521954 -7622 521986 -7386
rect 522222 -7622 522306 -7386
rect 522542 -7622 522574 -7386
rect 521954 -7654 522574 -7622
rect 531954 -6106 532574 14058
rect 534514 707718 535134 707750
rect 534514 707482 534546 707718
rect 534782 707482 534866 707718
rect 535102 707482 535134 707718
rect 534514 707398 535134 707482
rect 534514 707162 534546 707398
rect 534782 707162 534866 707398
rect 535102 707162 535134 707398
rect 534514 673174 535134 707162
rect 534514 672938 534546 673174
rect 534782 672938 534866 673174
rect 535102 672938 535134 673174
rect 534514 672854 535134 672938
rect 534514 672618 534546 672854
rect 534782 672618 534866 672854
rect 535102 672618 535134 672854
rect 534514 637174 535134 672618
rect 534514 636938 534546 637174
rect 534782 636938 534866 637174
rect 535102 636938 535134 637174
rect 534514 636854 535134 636938
rect 534514 636618 534546 636854
rect 534782 636618 534866 636854
rect 535102 636618 535134 636854
rect 534514 601174 535134 636618
rect 534514 600938 534546 601174
rect 534782 600938 534866 601174
rect 535102 600938 535134 601174
rect 534514 600854 535134 600938
rect 534514 600618 534546 600854
rect 534782 600618 534866 600854
rect 535102 600618 535134 600854
rect 534514 565174 535134 600618
rect 534514 564938 534546 565174
rect 534782 564938 534866 565174
rect 535102 564938 535134 565174
rect 534514 564854 535134 564938
rect 534514 564618 534546 564854
rect 534782 564618 534866 564854
rect 535102 564618 535134 564854
rect 534514 529174 535134 564618
rect 534514 528938 534546 529174
rect 534782 528938 534866 529174
rect 535102 528938 535134 529174
rect 534514 528854 535134 528938
rect 534514 528618 534546 528854
rect 534782 528618 534866 528854
rect 535102 528618 535134 528854
rect 534514 493174 535134 528618
rect 534514 492938 534546 493174
rect 534782 492938 534866 493174
rect 535102 492938 535134 493174
rect 534514 492854 535134 492938
rect 534514 492618 534546 492854
rect 534782 492618 534866 492854
rect 535102 492618 535134 492854
rect 534514 457174 535134 492618
rect 534514 456938 534546 457174
rect 534782 456938 534866 457174
rect 535102 456938 535134 457174
rect 534514 456854 535134 456938
rect 534514 456618 534546 456854
rect 534782 456618 534866 456854
rect 535102 456618 535134 456854
rect 534514 421174 535134 456618
rect 534514 420938 534546 421174
rect 534782 420938 534866 421174
rect 535102 420938 535134 421174
rect 534514 420854 535134 420938
rect 534514 420618 534546 420854
rect 534782 420618 534866 420854
rect 535102 420618 535134 420854
rect 534514 385174 535134 420618
rect 534514 384938 534546 385174
rect 534782 384938 534866 385174
rect 535102 384938 535134 385174
rect 534514 384854 535134 384938
rect 534514 384618 534546 384854
rect 534782 384618 534866 384854
rect 535102 384618 535134 384854
rect 534514 349174 535134 384618
rect 534514 348938 534546 349174
rect 534782 348938 534866 349174
rect 535102 348938 535134 349174
rect 534514 348854 535134 348938
rect 534514 348618 534546 348854
rect 534782 348618 534866 348854
rect 535102 348618 535134 348854
rect 534514 313174 535134 348618
rect 534514 312938 534546 313174
rect 534782 312938 534866 313174
rect 535102 312938 535134 313174
rect 534514 312854 535134 312938
rect 534514 312618 534546 312854
rect 534782 312618 534866 312854
rect 535102 312618 535134 312854
rect 534514 277174 535134 312618
rect 534514 276938 534546 277174
rect 534782 276938 534866 277174
rect 535102 276938 535134 277174
rect 534514 276854 535134 276938
rect 534514 276618 534546 276854
rect 534782 276618 534866 276854
rect 535102 276618 535134 276854
rect 534514 241174 535134 276618
rect 534514 240938 534546 241174
rect 534782 240938 534866 241174
rect 535102 240938 535134 241174
rect 534514 240854 535134 240938
rect 534514 240618 534546 240854
rect 534782 240618 534866 240854
rect 535102 240618 535134 240854
rect 534514 205174 535134 240618
rect 534514 204938 534546 205174
rect 534782 204938 534866 205174
rect 535102 204938 535134 205174
rect 534514 204854 535134 204938
rect 534514 204618 534546 204854
rect 534782 204618 534866 204854
rect 535102 204618 535134 204854
rect 534514 169174 535134 204618
rect 534514 168938 534546 169174
rect 534782 168938 534866 169174
rect 535102 168938 535134 169174
rect 534514 168854 535134 168938
rect 534514 168618 534546 168854
rect 534782 168618 534866 168854
rect 535102 168618 535134 168854
rect 534514 133174 535134 168618
rect 534514 132938 534546 133174
rect 534782 132938 534866 133174
rect 535102 132938 535134 133174
rect 534514 132854 535134 132938
rect 534514 132618 534546 132854
rect 534782 132618 534866 132854
rect 535102 132618 535134 132854
rect 534514 97174 535134 132618
rect 534514 96938 534546 97174
rect 534782 96938 534866 97174
rect 535102 96938 535134 97174
rect 534514 96854 535134 96938
rect 534514 96618 534546 96854
rect 534782 96618 534866 96854
rect 535102 96618 535134 96854
rect 534514 61174 535134 96618
rect 534514 60938 534546 61174
rect 534782 60938 534866 61174
rect 535102 60938 535134 61174
rect 534514 60854 535134 60938
rect 534514 60618 534546 60854
rect 534782 60618 534866 60854
rect 535102 60618 535134 60854
rect 534514 25174 535134 60618
rect 534514 24938 534546 25174
rect 534782 24938 534866 25174
rect 535102 24938 535134 25174
rect 534514 24854 535134 24938
rect 534514 24618 534546 24854
rect 534782 24618 534866 24854
rect 535102 24618 535134 24854
rect 534514 -3226 535134 24618
rect 534514 -3462 534546 -3226
rect 534782 -3462 534866 -3226
rect 535102 -3462 535134 -3226
rect 534514 -3546 535134 -3462
rect 534514 -3782 534546 -3546
rect 534782 -3782 534866 -3546
rect 535102 -3782 535134 -3546
rect 534514 -3814 535134 -3782
rect 538234 676894 538854 709082
rect 538234 676658 538266 676894
rect 538502 676658 538586 676894
rect 538822 676658 538854 676894
rect 538234 676574 538854 676658
rect 538234 676338 538266 676574
rect 538502 676338 538586 676574
rect 538822 676338 538854 676574
rect 538234 640894 538854 676338
rect 538234 640658 538266 640894
rect 538502 640658 538586 640894
rect 538822 640658 538854 640894
rect 538234 640574 538854 640658
rect 538234 640338 538266 640574
rect 538502 640338 538586 640574
rect 538822 640338 538854 640574
rect 538234 604894 538854 640338
rect 538234 604658 538266 604894
rect 538502 604658 538586 604894
rect 538822 604658 538854 604894
rect 538234 604574 538854 604658
rect 538234 604338 538266 604574
rect 538502 604338 538586 604574
rect 538822 604338 538854 604574
rect 538234 568894 538854 604338
rect 538234 568658 538266 568894
rect 538502 568658 538586 568894
rect 538822 568658 538854 568894
rect 538234 568574 538854 568658
rect 538234 568338 538266 568574
rect 538502 568338 538586 568574
rect 538822 568338 538854 568574
rect 538234 532894 538854 568338
rect 538234 532658 538266 532894
rect 538502 532658 538586 532894
rect 538822 532658 538854 532894
rect 538234 532574 538854 532658
rect 538234 532338 538266 532574
rect 538502 532338 538586 532574
rect 538822 532338 538854 532574
rect 538234 496894 538854 532338
rect 538234 496658 538266 496894
rect 538502 496658 538586 496894
rect 538822 496658 538854 496894
rect 538234 496574 538854 496658
rect 538234 496338 538266 496574
rect 538502 496338 538586 496574
rect 538822 496338 538854 496574
rect 538234 460894 538854 496338
rect 538234 460658 538266 460894
rect 538502 460658 538586 460894
rect 538822 460658 538854 460894
rect 538234 460574 538854 460658
rect 538234 460338 538266 460574
rect 538502 460338 538586 460574
rect 538822 460338 538854 460574
rect 538234 424894 538854 460338
rect 538234 424658 538266 424894
rect 538502 424658 538586 424894
rect 538822 424658 538854 424894
rect 538234 424574 538854 424658
rect 538234 424338 538266 424574
rect 538502 424338 538586 424574
rect 538822 424338 538854 424574
rect 538234 388894 538854 424338
rect 538234 388658 538266 388894
rect 538502 388658 538586 388894
rect 538822 388658 538854 388894
rect 538234 388574 538854 388658
rect 538234 388338 538266 388574
rect 538502 388338 538586 388574
rect 538822 388338 538854 388574
rect 538234 352894 538854 388338
rect 538234 352658 538266 352894
rect 538502 352658 538586 352894
rect 538822 352658 538854 352894
rect 538234 352574 538854 352658
rect 538234 352338 538266 352574
rect 538502 352338 538586 352574
rect 538822 352338 538854 352574
rect 538234 316894 538854 352338
rect 538234 316658 538266 316894
rect 538502 316658 538586 316894
rect 538822 316658 538854 316894
rect 538234 316574 538854 316658
rect 538234 316338 538266 316574
rect 538502 316338 538586 316574
rect 538822 316338 538854 316574
rect 538234 280894 538854 316338
rect 538234 280658 538266 280894
rect 538502 280658 538586 280894
rect 538822 280658 538854 280894
rect 538234 280574 538854 280658
rect 538234 280338 538266 280574
rect 538502 280338 538586 280574
rect 538822 280338 538854 280574
rect 538234 244894 538854 280338
rect 538234 244658 538266 244894
rect 538502 244658 538586 244894
rect 538822 244658 538854 244894
rect 538234 244574 538854 244658
rect 538234 244338 538266 244574
rect 538502 244338 538586 244574
rect 538822 244338 538854 244574
rect 538234 208894 538854 244338
rect 538234 208658 538266 208894
rect 538502 208658 538586 208894
rect 538822 208658 538854 208894
rect 538234 208574 538854 208658
rect 538234 208338 538266 208574
rect 538502 208338 538586 208574
rect 538822 208338 538854 208574
rect 538234 172894 538854 208338
rect 538234 172658 538266 172894
rect 538502 172658 538586 172894
rect 538822 172658 538854 172894
rect 538234 172574 538854 172658
rect 538234 172338 538266 172574
rect 538502 172338 538586 172574
rect 538822 172338 538854 172574
rect 538234 136894 538854 172338
rect 538234 136658 538266 136894
rect 538502 136658 538586 136894
rect 538822 136658 538854 136894
rect 538234 136574 538854 136658
rect 538234 136338 538266 136574
rect 538502 136338 538586 136574
rect 538822 136338 538854 136574
rect 538234 100894 538854 136338
rect 538234 100658 538266 100894
rect 538502 100658 538586 100894
rect 538822 100658 538854 100894
rect 538234 100574 538854 100658
rect 538234 100338 538266 100574
rect 538502 100338 538586 100574
rect 538822 100338 538854 100574
rect 538234 64894 538854 100338
rect 538234 64658 538266 64894
rect 538502 64658 538586 64894
rect 538822 64658 538854 64894
rect 538234 64574 538854 64658
rect 538234 64338 538266 64574
rect 538502 64338 538586 64574
rect 538822 64338 538854 64574
rect 538234 28894 538854 64338
rect 538234 28658 538266 28894
rect 538502 28658 538586 28894
rect 538822 28658 538854 28894
rect 538234 28574 538854 28658
rect 538234 28338 538266 28574
rect 538502 28338 538586 28574
rect 538822 28338 538854 28574
rect 538234 -5146 538854 28338
rect 540794 704838 541414 705830
rect 540794 704602 540826 704838
rect 541062 704602 541146 704838
rect 541382 704602 541414 704838
rect 540794 704518 541414 704602
rect 540794 704282 540826 704518
rect 541062 704282 541146 704518
rect 541382 704282 541414 704518
rect 540794 687454 541414 704282
rect 540794 687218 540826 687454
rect 541062 687218 541146 687454
rect 541382 687218 541414 687454
rect 540794 687134 541414 687218
rect 540794 686898 540826 687134
rect 541062 686898 541146 687134
rect 541382 686898 541414 687134
rect 540794 651454 541414 686898
rect 540794 651218 540826 651454
rect 541062 651218 541146 651454
rect 541382 651218 541414 651454
rect 540794 651134 541414 651218
rect 540794 650898 540826 651134
rect 541062 650898 541146 651134
rect 541382 650898 541414 651134
rect 540794 615454 541414 650898
rect 540794 615218 540826 615454
rect 541062 615218 541146 615454
rect 541382 615218 541414 615454
rect 540794 615134 541414 615218
rect 540794 614898 540826 615134
rect 541062 614898 541146 615134
rect 541382 614898 541414 615134
rect 540794 579454 541414 614898
rect 540794 579218 540826 579454
rect 541062 579218 541146 579454
rect 541382 579218 541414 579454
rect 540794 579134 541414 579218
rect 540794 578898 540826 579134
rect 541062 578898 541146 579134
rect 541382 578898 541414 579134
rect 540794 543454 541414 578898
rect 540794 543218 540826 543454
rect 541062 543218 541146 543454
rect 541382 543218 541414 543454
rect 540794 543134 541414 543218
rect 540794 542898 540826 543134
rect 541062 542898 541146 543134
rect 541382 542898 541414 543134
rect 540794 507454 541414 542898
rect 540794 507218 540826 507454
rect 541062 507218 541146 507454
rect 541382 507218 541414 507454
rect 540794 507134 541414 507218
rect 540794 506898 540826 507134
rect 541062 506898 541146 507134
rect 541382 506898 541414 507134
rect 540794 471454 541414 506898
rect 540794 471218 540826 471454
rect 541062 471218 541146 471454
rect 541382 471218 541414 471454
rect 540794 471134 541414 471218
rect 540794 470898 540826 471134
rect 541062 470898 541146 471134
rect 541382 470898 541414 471134
rect 540794 435454 541414 470898
rect 540794 435218 540826 435454
rect 541062 435218 541146 435454
rect 541382 435218 541414 435454
rect 540794 435134 541414 435218
rect 540794 434898 540826 435134
rect 541062 434898 541146 435134
rect 541382 434898 541414 435134
rect 540794 399454 541414 434898
rect 540794 399218 540826 399454
rect 541062 399218 541146 399454
rect 541382 399218 541414 399454
rect 540794 399134 541414 399218
rect 540794 398898 540826 399134
rect 541062 398898 541146 399134
rect 541382 398898 541414 399134
rect 540794 363454 541414 398898
rect 540794 363218 540826 363454
rect 541062 363218 541146 363454
rect 541382 363218 541414 363454
rect 540794 363134 541414 363218
rect 540794 362898 540826 363134
rect 541062 362898 541146 363134
rect 541382 362898 541414 363134
rect 540794 327454 541414 362898
rect 540794 327218 540826 327454
rect 541062 327218 541146 327454
rect 541382 327218 541414 327454
rect 540794 327134 541414 327218
rect 540794 326898 540826 327134
rect 541062 326898 541146 327134
rect 541382 326898 541414 327134
rect 540794 291454 541414 326898
rect 540794 291218 540826 291454
rect 541062 291218 541146 291454
rect 541382 291218 541414 291454
rect 540794 291134 541414 291218
rect 540794 290898 540826 291134
rect 541062 290898 541146 291134
rect 541382 290898 541414 291134
rect 540794 255454 541414 290898
rect 540794 255218 540826 255454
rect 541062 255218 541146 255454
rect 541382 255218 541414 255454
rect 540794 255134 541414 255218
rect 540794 254898 540826 255134
rect 541062 254898 541146 255134
rect 541382 254898 541414 255134
rect 540794 219454 541414 254898
rect 540794 219218 540826 219454
rect 541062 219218 541146 219454
rect 541382 219218 541414 219454
rect 540794 219134 541414 219218
rect 540794 218898 540826 219134
rect 541062 218898 541146 219134
rect 541382 218898 541414 219134
rect 540794 183454 541414 218898
rect 540794 183218 540826 183454
rect 541062 183218 541146 183454
rect 541382 183218 541414 183454
rect 540794 183134 541414 183218
rect 540794 182898 540826 183134
rect 541062 182898 541146 183134
rect 541382 182898 541414 183134
rect 540794 147454 541414 182898
rect 540794 147218 540826 147454
rect 541062 147218 541146 147454
rect 541382 147218 541414 147454
rect 540794 147134 541414 147218
rect 540794 146898 540826 147134
rect 541062 146898 541146 147134
rect 541382 146898 541414 147134
rect 540794 111454 541414 146898
rect 540794 111218 540826 111454
rect 541062 111218 541146 111454
rect 541382 111218 541414 111454
rect 540794 111134 541414 111218
rect 540794 110898 540826 111134
rect 541062 110898 541146 111134
rect 541382 110898 541414 111134
rect 540794 75454 541414 110898
rect 540794 75218 540826 75454
rect 541062 75218 541146 75454
rect 541382 75218 541414 75454
rect 540794 75134 541414 75218
rect 540794 74898 540826 75134
rect 541062 74898 541146 75134
rect 541382 74898 541414 75134
rect 540794 39454 541414 74898
rect 540794 39218 540826 39454
rect 541062 39218 541146 39454
rect 541382 39218 541414 39454
rect 540794 39134 541414 39218
rect 540794 38898 540826 39134
rect 541062 38898 541146 39134
rect 541382 38898 541414 39134
rect 540794 3454 541414 38898
rect 540794 3218 540826 3454
rect 541062 3218 541146 3454
rect 541382 3218 541414 3454
rect 540794 3134 541414 3218
rect 540794 2898 540826 3134
rect 541062 2898 541146 3134
rect 541382 2898 541414 3134
rect 540794 -346 541414 2898
rect 540794 -582 540826 -346
rect 541062 -582 541146 -346
rect 541382 -582 541414 -346
rect 540794 -666 541414 -582
rect 540794 -902 540826 -666
rect 541062 -902 541146 -666
rect 541382 -902 541414 -666
rect 540794 -1894 541414 -902
rect 541954 680614 542574 711002
rect 551954 710598 552574 711590
rect 551954 710362 551986 710598
rect 552222 710362 552306 710598
rect 552542 710362 552574 710598
rect 551954 710278 552574 710362
rect 551954 710042 551986 710278
rect 552222 710042 552306 710278
rect 552542 710042 552574 710278
rect 548234 708678 548854 709670
rect 548234 708442 548266 708678
rect 548502 708442 548586 708678
rect 548822 708442 548854 708678
rect 548234 708358 548854 708442
rect 548234 708122 548266 708358
rect 548502 708122 548586 708358
rect 548822 708122 548854 708358
rect 541954 680378 541986 680614
rect 542222 680378 542306 680614
rect 542542 680378 542574 680614
rect 541954 680294 542574 680378
rect 541954 680058 541986 680294
rect 542222 680058 542306 680294
rect 542542 680058 542574 680294
rect 541954 644614 542574 680058
rect 541954 644378 541986 644614
rect 542222 644378 542306 644614
rect 542542 644378 542574 644614
rect 541954 644294 542574 644378
rect 541954 644058 541986 644294
rect 542222 644058 542306 644294
rect 542542 644058 542574 644294
rect 541954 608614 542574 644058
rect 541954 608378 541986 608614
rect 542222 608378 542306 608614
rect 542542 608378 542574 608614
rect 541954 608294 542574 608378
rect 541954 608058 541986 608294
rect 542222 608058 542306 608294
rect 542542 608058 542574 608294
rect 541954 572614 542574 608058
rect 541954 572378 541986 572614
rect 542222 572378 542306 572614
rect 542542 572378 542574 572614
rect 541954 572294 542574 572378
rect 541954 572058 541986 572294
rect 542222 572058 542306 572294
rect 542542 572058 542574 572294
rect 541954 536614 542574 572058
rect 541954 536378 541986 536614
rect 542222 536378 542306 536614
rect 542542 536378 542574 536614
rect 541954 536294 542574 536378
rect 541954 536058 541986 536294
rect 542222 536058 542306 536294
rect 542542 536058 542574 536294
rect 541954 500614 542574 536058
rect 541954 500378 541986 500614
rect 542222 500378 542306 500614
rect 542542 500378 542574 500614
rect 541954 500294 542574 500378
rect 541954 500058 541986 500294
rect 542222 500058 542306 500294
rect 542542 500058 542574 500294
rect 541954 464614 542574 500058
rect 541954 464378 541986 464614
rect 542222 464378 542306 464614
rect 542542 464378 542574 464614
rect 541954 464294 542574 464378
rect 541954 464058 541986 464294
rect 542222 464058 542306 464294
rect 542542 464058 542574 464294
rect 541954 428614 542574 464058
rect 541954 428378 541986 428614
rect 542222 428378 542306 428614
rect 542542 428378 542574 428614
rect 541954 428294 542574 428378
rect 541954 428058 541986 428294
rect 542222 428058 542306 428294
rect 542542 428058 542574 428294
rect 541954 392614 542574 428058
rect 541954 392378 541986 392614
rect 542222 392378 542306 392614
rect 542542 392378 542574 392614
rect 541954 392294 542574 392378
rect 541954 392058 541986 392294
rect 542222 392058 542306 392294
rect 542542 392058 542574 392294
rect 541954 356614 542574 392058
rect 541954 356378 541986 356614
rect 542222 356378 542306 356614
rect 542542 356378 542574 356614
rect 541954 356294 542574 356378
rect 541954 356058 541986 356294
rect 542222 356058 542306 356294
rect 542542 356058 542574 356294
rect 541954 320614 542574 356058
rect 541954 320378 541986 320614
rect 542222 320378 542306 320614
rect 542542 320378 542574 320614
rect 541954 320294 542574 320378
rect 541954 320058 541986 320294
rect 542222 320058 542306 320294
rect 542542 320058 542574 320294
rect 541954 284614 542574 320058
rect 541954 284378 541986 284614
rect 542222 284378 542306 284614
rect 542542 284378 542574 284614
rect 541954 284294 542574 284378
rect 541954 284058 541986 284294
rect 542222 284058 542306 284294
rect 542542 284058 542574 284294
rect 541954 248614 542574 284058
rect 541954 248378 541986 248614
rect 542222 248378 542306 248614
rect 542542 248378 542574 248614
rect 541954 248294 542574 248378
rect 541954 248058 541986 248294
rect 542222 248058 542306 248294
rect 542542 248058 542574 248294
rect 541954 212614 542574 248058
rect 541954 212378 541986 212614
rect 542222 212378 542306 212614
rect 542542 212378 542574 212614
rect 541954 212294 542574 212378
rect 541954 212058 541986 212294
rect 542222 212058 542306 212294
rect 542542 212058 542574 212294
rect 541954 176614 542574 212058
rect 541954 176378 541986 176614
rect 542222 176378 542306 176614
rect 542542 176378 542574 176614
rect 541954 176294 542574 176378
rect 541954 176058 541986 176294
rect 542222 176058 542306 176294
rect 542542 176058 542574 176294
rect 541954 140614 542574 176058
rect 541954 140378 541986 140614
rect 542222 140378 542306 140614
rect 542542 140378 542574 140614
rect 541954 140294 542574 140378
rect 541954 140058 541986 140294
rect 542222 140058 542306 140294
rect 542542 140058 542574 140294
rect 541954 104614 542574 140058
rect 541954 104378 541986 104614
rect 542222 104378 542306 104614
rect 542542 104378 542574 104614
rect 541954 104294 542574 104378
rect 541954 104058 541986 104294
rect 542222 104058 542306 104294
rect 542542 104058 542574 104294
rect 541954 68614 542574 104058
rect 541954 68378 541986 68614
rect 542222 68378 542306 68614
rect 542542 68378 542574 68614
rect 541954 68294 542574 68378
rect 541954 68058 541986 68294
rect 542222 68058 542306 68294
rect 542542 68058 542574 68294
rect 541954 32614 542574 68058
rect 541954 32378 541986 32614
rect 542222 32378 542306 32614
rect 542542 32378 542574 32614
rect 541954 32294 542574 32378
rect 541954 32058 541986 32294
rect 542222 32058 542306 32294
rect 542542 32058 542574 32294
rect 538234 -5382 538266 -5146
rect 538502 -5382 538586 -5146
rect 538822 -5382 538854 -5146
rect 538234 -5466 538854 -5382
rect 538234 -5702 538266 -5466
rect 538502 -5702 538586 -5466
rect 538822 -5702 538854 -5466
rect 538234 -5734 538854 -5702
rect 531954 -6342 531986 -6106
rect 532222 -6342 532306 -6106
rect 532542 -6342 532574 -6106
rect 531954 -6426 532574 -6342
rect 531954 -6662 531986 -6426
rect 532222 -6662 532306 -6426
rect 532542 -6662 532574 -6426
rect 531954 -7654 532574 -6662
rect 541954 -7066 542574 32058
rect 544514 706758 545134 707750
rect 544514 706522 544546 706758
rect 544782 706522 544866 706758
rect 545102 706522 545134 706758
rect 544514 706438 545134 706522
rect 544514 706202 544546 706438
rect 544782 706202 544866 706438
rect 545102 706202 545134 706438
rect 544514 691174 545134 706202
rect 544514 690938 544546 691174
rect 544782 690938 544866 691174
rect 545102 690938 545134 691174
rect 544514 690854 545134 690938
rect 544514 690618 544546 690854
rect 544782 690618 544866 690854
rect 545102 690618 545134 690854
rect 544514 655174 545134 690618
rect 544514 654938 544546 655174
rect 544782 654938 544866 655174
rect 545102 654938 545134 655174
rect 544514 654854 545134 654938
rect 544514 654618 544546 654854
rect 544782 654618 544866 654854
rect 545102 654618 545134 654854
rect 544514 619174 545134 654618
rect 544514 618938 544546 619174
rect 544782 618938 544866 619174
rect 545102 618938 545134 619174
rect 544514 618854 545134 618938
rect 544514 618618 544546 618854
rect 544782 618618 544866 618854
rect 545102 618618 545134 618854
rect 544514 583174 545134 618618
rect 544514 582938 544546 583174
rect 544782 582938 544866 583174
rect 545102 582938 545134 583174
rect 544514 582854 545134 582938
rect 544514 582618 544546 582854
rect 544782 582618 544866 582854
rect 545102 582618 545134 582854
rect 544514 547174 545134 582618
rect 544514 546938 544546 547174
rect 544782 546938 544866 547174
rect 545102 546938 545134 547174
rect 544514 546854 545134 546938
rect 544514 546618 544546 546854
rect 544782 546618 544866 546854
rect 545102 546618 545134 546854
rect 544514 511174 545134 546618
rect 544514 510938 544546 511174
rect 544782 510938 544866 511174
rect 545102 510938 545134 511174
rect 544514 510854 545134 510938
rect 544514 510618 544546 510854
rect 544782 510618 544866 510854
rect 545102 510618 545134 510854
rect 544514 475174 545134 510618
rect 544514 474938 544546 475174
rect 544782 474938 544866 475174
rect 545102 474938 545134 475174
rect 544514 474854 545134 474938
rect 544514 474618 544546 474854
rect 544782 474618 544866 474854
rect 545102 474618 545134 474854
rect 544514 439174 545134 474618
rect 544514 438938 544546 439174
rect 544782 438938 544866 439174
rect 545102 438938 545134 439174
rect 544514 438854 545134 438938
rect 544514 438618 544546 438854
rect 544782 438618 544866 438854
rect 545102 438618 545134 438854
rect 544514 403174 545134 438618
rect 544514 402938 544546 403174
rect 544782 402938 544866 403174
rect 545102 402938 545134 403174
rect 544514 402854 545134 402938
rect 544514 402618 544546 402854
rect 544782 402618 544866 402854
rect 545102 402618 545134 402854
rect 544514 367174 545134 402618
rect 544514 366938 544546 367174
rect 544782 366938 544866 367174
rect 545102 366938 545134 367174
rect 544514 366854 545134 366938
rect 544514 366618 544546 366854
rect 544782 366618 544866 366854
rect 545102 366618 545134 366854
rect 544514 331174 545134 366618
rect 544514 330938 544546 331174
rect 544782 330938 544866 331174
rect 545102 330938 545134 331174
rect 544514 330854 545134 330938
rect 544514 330618 544546 330854
rect 544782 330618 544866 330854
rect 545102 330618 545134 330854
rect 544514 295174 545134 330618
rect 544514 294938 544546 295174
rect 544782 294938 544866 295174
rect 545102 294938 545134 295174
rect 544514 294854 545134 294938
rect 544514 294618 544546 294854
rect 544782 294618 544866 294854
rect 545102 294618 545134 294854
rect 544514 259174 545134 294618
rect 544514 258938 544546 259174
rect 544782 258938 544866 259174
rect 545102 258938 545134 259174
rect 544514 258854 545134 258938
rect 544514 258618 544546 258854
rect 544782 258618 544866 258854
rect 545102 258618 545134 258854
rect 544514 223174 545134 258618
rect 544514 222938 544546 223174
rect 544782 222938 544866 223174
rect 545102 222938 545134 223174
rect 544514 222854 545134 222938
rect 544514 222618 544546 222854
rect 544782 222618 544866 222854
rect 545102 222618 545134 222854
rect 544514 187174 545134 222618
rect 544514 186938 544546 187174
rect 544782 186938 544866 187174
rect 545102 186938 545134 187174
rect 544514 186854 545134 186938
rect 544514 186618 544546 186854
rect 544782 186618 544866 186854
rect 545102 186618 545134 186854
rect 544514 151174 545134 186618
rect 544514 150938 544546 151174
rect 544782 150938 544866 151174
rect 545102 150938 545134 151174
rect 544514 150854 545134 150938
rect 544514 150618 544546 150854
rect 544782 150618 544866 150854
rect 545102 150618 545134 150854
rect 544514 115174 545134 150618
rect 544514 114938 544546 115174
rect 544782 114938 544866 115174
rect 545102 114938 545134 115174
rect 544514 114854 545134 114938
rect 544514 114618 544546 114854
rect 544782 114618 544866 114854
rect 545102 114618 545134 114854
rect 544514 79174 545134 114618
rect 544514 78938 544546 79174
rect 544782 78938 544866 79174
rect 545102 78938 545134 79174
rect 544514 78854 545134 78938
rect 544514 78618 544546 78854
rect 544782 78618 544866 78854
rect 545102 78618 545134 78854
rect 544514 43174 545134 78618
rect 544514 42938 544546 43174
rect 544782 42938 544866 43174
rect 545102 42938 545134 43174
rect 544514 42854 545134 42938
rect 544514 42618 544546 42854
rect 544782 42618 544866 42854
rect 545102 42618 545134 42854
rect 544514 7174 545134 42618
rect 544514 6938 544546 7174
rect 544782 6938 544866 7174
rect 545102 6938 545134 7174
rect 544514 6854 545134 6938
rect 544514 6618 544546 6854
rect 544782 6618 544866 6854
rect 545102 6618 545134 6854
rect 544514 -2266 545134 6618
rect 544514 -2502 544546 -2266
rect 544782 -2502 544866 -2266
rect 545102 -2502 545134 -2266
rect 544514 -2586 545134 -2502
rect 544514 -2822 544546 -2586
rect 544782 -2822 544866 -2586
rect 545102 -2822 545134 -2586
rect 544514 -3814 545134 -2822
rect 548234 694894 548854 708122
rect 548234 694658 548266 694894
rect 548502 694658 548586 694894
rect 548822 694658 548854 694894
rect 548234 694574 548854 694658
rect 548234 694338 548266 694574
rect 548502 694338 548586 694574
rect 548822 694338 548854 694574
rect 548234 658894 548854 694338
rect 548234 658658 548266 658894
rect 548502 658658 548586 658894
rect 548822 658658 548854 658894
rect 548234 658574 548854 658658
rect 548234 658338 548266 658574
rect 548502 658338 548586 658574
rect 548822 658338 548854 658574
rect 548234 622894 548854 658338
rect 548234 622658 548266 622894
rect 548502 622658 548586 622894
rect 548822 622658 548854 622894
rect 548234 622574 548854 622658
rect 548234 622338 548266 622574
rect 548502 622338 548586 622574
rect 548822 622338 548854 622574
rect 548234 586894 548854 622338
rect 548234 586658 548266 586894
rect 548502 586658 548586 586894
rect 548822 586658 548854 586894
rect 548234 586574 548854 586658
rect 548234 586338 548266 586574
rect 548502 586338 548586 586574
rect 548822 586338 548854 586574
rect 548234 550894 548854 586338
rect 548234 550658 548266 550894
rect 548502 550658 548586 550894
rect 548822 550658 548854 550894
rect 548234 550574 548854 550658
rect 548234 550338 548266 550574
rect 548502 550338 548586 550574
rect 548822 550338 548854 550574
rect 548234 514894 548854 550338
rect 548234 514658 548266 514894
rect 548502 514658 548586 514894
rect 548822 514658 548854 514894
rect 548234 514574 548854 514658
rect 548234 514338 548266 514574
rect 548502 514338 548586 514574
rect 548822 514338 548854 514574
rect 548234 478894 548854 514338
rect 548234 478658 548266 478894
rect 548502 478658 548586 478894
rect 548822 478658 548854 478894
rect 548234 478574 548854 478658
rect 548234 478338 548266 478574
rect 548502 478338 548586 478574
rect 548822 478338 548854 478574
rect 548234 442894 548854 478338
rect 548234 442658 548266 442894
rect 548502 442658 548586 442894
rect 548822 442658 548854 442894
rect 548234 442574 548854 442658
rect 548234 442338 548266 442574
rect 548502 442338 548586 442574
rect 548822 442338 548854 442574
rect 548234 406894 548854 442338
rect 548234 406658 548266 406894
rect 548502 406658 548586 406894
rect 548822 406658 548854 406894
rect 548234 406574 548854 406658
rect 548234 406338 548266 406574
rect 548502 406338 548586 406574
rect 548822 406338 548854 406574
rect 548234 370894 548854 406338
rect 548234 370658 548266 370894
rect 548502 370658 548586 370894
rect 548822 370658 548854 370894
rect 548234 370574 548854 370658
rect 548234 370338 548266 370574
rect 548502 370338 548586 370574
rect 548822 370338 548854 370574
rect 548234 334894 548854 370338
rect 548234 334658 548266 334894
rect 548502 334658 548586 334894
rect 548822 334658 548854 334894
rect 548234 334574 548854 334658
rect 548234 334338 548266 334574
rect 548502 334338 548586 334574
rect 548822 334338 548854 334574
rect 548234 298894 548854 334338
rect 548234 298658 548266 298894
rect 548502 298658 548586 298894
rect 548822 298658 548854 298894
rect 548234 298574 548854 298658
rect 548234 298338 548266 298574
rect 548502 298338 548586 298574
rect 548822 298338 548854 298574
rect 548234 262894 548854 298338
rect 548234 262658 548266 262894
rect 548502 262658 548586 262894
rect 548822 262658 548854 262894
rect 548234 262574 548854 262658
rect 548234 262338 548266 262574
rect 548502 262338 548586 262574
rect 548822 262338 548854 262574
rect 548234 226894 548854 262338
rect 548234 226658 548266 226894
rect 548502 226658 548586 226894
rect 548822 226658 548854 226894
rect 548234 226574 548854 226658
rect 548234 226338 548266 226574
rect 548502 226338 548586 226574
rect 548822 226338 548854 226574
rect 548234 190894 548854 226338
rect 548234 190658 548266 190894
rect 548502 190658 548586 190894
rect 548822 190658 548854 190894
rect 548234 190574 548854 190658
rect 548234 190338 548266 190574
rect 548502 190338 548586 190574
rect 548822 190338 548854 190574
rect 548234 154894 548854 190338
rect 548234 154658 548266 154894
rect 548502 154658 548586 154894
rect 548822 154658 548854 154894
rect 548234 154574 548854 154658
rect 548234 154338 548266 154574
rect 548502 154338 548586 154574
rect 548822 154338 548854 154574
rect 548234 118894 548854 154338
rect 548234 118658 548266 118894
rect 548502 118658 548586 118894
rect 548822 118658 548854 118894
rect 548234 118574 548854 118658
rect 548234 118338 548266 118574
rect 548502 118338 548586 118574
rect 548822 118338 548854 118574
rect 548234 82894 548854 118338
rect 548234 82658 548266 82894
rect 548502 82658 548586 82894
rect 548822 82658 548854 82894
rect 548234 82574 548854 82658
rect 548234 82338 548266 82574
rect 548502 82338 548586 82574
rect 548822 82338 548854 82574
rect 548234 46894 548854 82338
rect 548234 46658 548266 46894
rect 548502 46658 548586 46894
rect 548822 46658 548854 46894
rect 548234 46574 548854 46658
rect 548234 46338 548266 46574
rect 548502 46338 548586 46574
rect 548822 46338 548854 46574
rect 548234 10894 548854 46338
rect 548234 10658 548266 10894
rect 548502 10658 548586 10894
rect 548822 10658 548854 10894
rect 548234 10574 548854 10658
rect 548234 10338 548266 10574
rect 548502 10338 548586 10574
rect 548822 10338 548854 10574
rect 548234 -4186 548854 10338
rect 550794 705798 551414 705830
rect 550794 705562 550826 705798
rect 551062 705562 551146 705798
rect 551382 705562 551414 705798
rect 550794 705478 551414 705562
rect 550794 705242 550826 705478
rect 551062 705242 551146 705478
rect 551382 705242 551414 705478
rect 550794 669454 551414 705242
rect 550794 669218 550826 669454
rect 551062 669218 551146 669454
rect 551382 669218 551414 669454
rect 550794 669134 551414 669218
rect 550794 668898 550826 669134
rect 551062 668898 551146 669134
rect 551382 668898 551414 669134
rect 550794 633454 551414 668898
rect 550794 633218 550826 633454
rect 551062 633218 551146 633454
rect 551382 633218 551414 633454
rect 550794 633134 551414 633218
rect 550794 632898 550826 633134
rect 551062 632898 551146 633134
rect 551382 632898 551414 633134
rect 550794 597454 551414 632898
rect 550794 597218 550826 597454
rect 551062 597218 551146 597454
rect 551382 597218 551414 597454
rect 550794 597134 551414 597218
rect 550794 596898 550826 597134
rect 551062 596898 551146 597134
rect 551382 596898 551414 597134
rect 550794 561454 551414 596898
rect 550794 561218 550826 561454
rect 551062 561218 551146 561454
rect 551382 561218 551414 561454
rect 550794 561134 551414 561218
rect 550794 560898 550826 561134
rect 551062 560898 551146 561134
rect 551382 560898 551414 561134
rect 550794 525454 551414 560898
rect 550794 525218 550826 525454
rect 551062 525218 551146 525454
rect 551382 525218 551414 525454
rect 550794 525134 551414 525218
rect 550794 524898 550826 525134
rect 551062 524898 551146 525134
rect 551382 524898 551414 525134
rect 550794 489454 551414 524898
rect 550794 489218 550826 489454
rect 551062 489218 551146 489454
rect 551382 489218 551414 489454
rect 550794 489134 551414 489218
rect 550794 488898 550826 489134
rect 551062 488898 551146 489134
rect 551382 488898 551414 489134
rect 550794 453454 551414 488898
rect 550794 453218 550826 453454
rect 551062 453218 551146 453454
rect 551382 453218 551414 453454
rect 550794 453134 551414 453218
rect 550794 452898 550826 453134
rect 551062 452898 551146 453134
rect 551382 452898 551414 453134
rect 550794 417454 551414 452898
rect 550794 417218 550826 417454
rect 551062 417218 551146 417454
rect 551382 417218 551414 417454
rect 550794 417134 551414 417218
rect 550794 416898 550826 417134
rect 551062 416898 551146 417134
rect 551382 416898 551414 417134
rect 550794 381454 551414 416898
rect 550794 381218 550826 381454
rect 551062 381218 551146 381454
rect 551382 381218 551414 381454
rect 550794 381134 551414 381218
rect 550794 380898 550826 381134
rect 551062 380898 551146 381134
rect 551382 380898 551414 381134
rect 550794 345454 551414 380898
rect 550794 345218 550826 345454
rect 551062 345218 551146 345454
rect 551382 345218 551414 345454
rect 550794 345134 551414 345218
rect 550794 344898 550826 345134
rect 551062 344898 551146 345134
rect 551382 344898 551414 345134
rect 550794 309454 551414 344898
rect 550794 309218 550826 309454
rect 551062 309218 551146 309454
rect 551382 309218 551414 309454
rect 550794 309134 551414 309218
rect 550794 308898 550826 309134
rect 551062 308898 551146 309134
rect 551382 308898 551414 309134
rect 550794 273454 551414 308898
rect 550794 273218 550826 273454
rect 551062 273218 551146 273454
rect 551382 273218 551414 273454
rect 550794 273134 551414 273218
rect 550794 272898 550826 273134
rect 551062 272898 551146 273134
rect 551382 272898 551414 273134
rect 550794 237454 551414 272898
rect 550794 237218 550826 237454
rect 551062 237218 551146 237454
rect 551382 237218 551414 237454
rect 550794 237134 551414 237218
rect 550794 236898 550826 237134
rect 551062 236898 551146 237134
rect 551382 236898 551414 237134
rect 550794 201454 551414 236898
rect 550794 201218 550826 201454
rect 551062 201218 551146 201454
rect 551382 201218 551414 201454
rect 550794 201134 551414 201218
rect 550794 200898 550826 201134
rect 551062 200898 551146 201134
rect 551382 200898 551414 201134
rect 550794 165454 551414 200898
rect 550794 165218 550826 165454
rect 551062 165218 551146 165454
rect 551382 165218 551414 165454
rect 550794 165134 551414 165218
rect 550794 164898 550826 165134
rect 551062 164898 551146 165134
rect 551382 164898 551414 165134
rect 550794 129454 551414 164898
rect 550794 129218 550826 129454
rect 551062 129218 551146 129454
rect 551382 129218 551414 129454
rect 550794 129134 551414 129218
rect 550794 128898 550826 129134
rect 551062 128898 551146 129134
rect 551382 128898 551414 129134
rect 550794 93454 551414 128898
rect 550794 93218 550826 93454
rect 551062 93218 551146 93454
rect 551382 93218 551414 93454
rect 550794 93134 551414 93218
rect 550794 92898 550826 93134
rect 551062 92898 551146 93134
rect 551382 92898 551414 93134
rect 550794 57454 551414 92898
rect 550794 57218 550826 57454
rect 551062 57218 551146 57454
rect 551382 57218 551414 57454
rect 550794 57134 551414 57218
rect 550794 56898 550826 57134
rect 551062 56898 551146 57134
rect 551382 56898 551414 57134
rect 550794 21454 551414 56898
rect 550794 21218 550826 21454
rect 551062 21218 551146 21454
rect 551382 21218 551414 21454
rect 550794 21134 551414 21218
rect 550794 20898 550826 21134
rect 551062 20898 551146 21134
rect 551382 20898 551414 21134
rect 550794 -1306 551414 20898
rect 550794 -1542 550826 -1306
rect 551062 -1542 551146 -1306
rect 551382 -1542 551414 -1306
rect 550794 -1626 551414 -1542
rect 550794 -1862 550826 -1626
rect 551062 -1862 551146 -1626
rect 551382 -1862 551414 -1626
rect 550794 -1894 551414 -1862
rect 551954 698614 552574 710042
rect 561954 711558 562574 711590
rect 561954 711322 561986 711558
rect 562222 711322 562306 711558
rect 562542 711322 562574 711558
rect 561954 711238 562574 711322
rect 561954 711002 561986 711238
rect 562222 711002 562306 711238
rect 562542 711002 562574 711238
rect 558234 709638 558854 709670
rect 558234 709402 558266 709638
rect 558502 709402 558586 709638
rect 558822 709402 558854 709638
rect 558234 709318 558854 709402
rect 558234 709082 558266 709318
rect 558502 709082 558586 709318
rect 558822 709082 558854 709318
rect 551954 698378 551986 698614
rect 552222 698378 552306 698614
rect 552542 698378 552574 698614
rect 551954 698294 552574 698378
rect 551954 698058 551986 698294
rect 552222 698058 552306 698294
rect 552542 698058 552574 698294
rect 551954 662614 552574 698058
rect 551954 662378 551986 662614
rect 552222 662378 552306 662614
rect 552542 662378 552574 662614
rect 551954 662294 552574 662378
rect 551954 662058 551986 662294
rect 552222 662058 552306 662294
rect 552542 662058 552574 662294
rect 551954 626614 552574 662058
rect 551954 626378 551986 626614
rect 552222 626378 552306 626614
rect 552542 626378 552574 626614
rect 551954 626294 552574 626378
rect 551954 626058 551986 626294
rect 552222 626058 552306 626294
rect 552542 626058 552574 626294
rect 551954 590614 552574 626058
rect 551954 590378 551986 590614
rect 552222 590378 552306 590614
rect 552542 590378 552574 590614
rect 551954 590294 552574 590378
rect 551954 590058 551986 590294
rect 552222 590058 552306 590294
rect 552542 590058 552574 590294
rect 551954 554614 552574 590058
rect 551954 554378 551986 554614
rect 552222 554378 552306 554614
rect 552542 554378 552574 554614
rect 551954 554294 552574 554378
rect 551954 554058 551986 554294
rect 552222 554058 552306 554294
rect 552542 554058 552574 554294
rect 551954 518614 552574 554058
rect 551954 518378 551986 518614
rect 552222 518378 552306 518614
rect 552542 518378 552574 518614
rect 551954 518294 552574 518378
rect 551954 518058 551986 518294
rect 552222 518058 552306 518294
rect 552542 518058 552574 518294
rect 551954 482614 552574 518058
rect 551954 482378 551986 482614
rect 552222 482378 552306 482614
rect 552542 482378 552574 482614
rect 551954 482294 552574 482378
rect 551954 482058 551986 482294
rect 552222 482058 552306 482294
rect 552542 482058 552574 482294
rect 551954 446614 552574 482058
rect 551954 446378 551986 446614
rect 552222 446378 552306 446614
rect 552542 446378 552574 446614
rect 551954 446294 552574 446378
rect 551954 446058 551986 446294
rect 552222 446058 552306 446294
rect 552542 446058 552574 446294
rect 551954 410614 552574 446058
rect 551954 410378 551986 410614
rect 552222 410378 552306 410614
rect 552542 410378 552574 410614
rect 551954 410294 552574 410378
rect 551954 410058 551986 410294
rect 552222 410058 552306 410294
rect 552542 410058 552574 410294
rect 551954 374614 552574 410058
rect 551954 374378 551986 374614
rect 552222 374378 552306 374614
rect 552542 374378 552574 374614
rect 551954 374294 552574 374378
rect 551954 374058 551986 374294
rect 552222 374058 552306 374294
rect 552542 374058 552574 374294
rect 551954 338614 552574 374058
rect 551954 338378 551986 338614
rect 552222 338378 552306 338614
rect 552542 338378 552574 338614
rect 551954 338294 552574 338378
rect 551954 338058 551986 338294
rect 552222 338058 552306 338294
rect 552542 338058 552574 338294
rect 551954 302614 552574 338058
rect 551954 302378 551986 302614
rect 552222 302378 552306 302614
rect 552542 302378 552574 302614
rect 551954 302294 552574 302378
rect 551954 302058 551986 302294
rect 552222 302058 552306 302294
rect 552542 302058 552574 302294
rect 551954 266614 552574 302058
rect 551954 266378 551986 266614
rect 552222 266378 552306 266614
rect 552542 266378 552574 266614
rect 551954 266294 552574 266378
rect 551954 266058 551986 266294
rect 552222 266058 552306 266294
rect 552542 266058 552574 266294
rect 551954 230614 552574 266058
rect 551954 230378 551986 230614
rect 552222 230378 552306 230614
rect 552542 230378 552574 230614
rect 551954 230294 552574 230378
rect 551954 230058 551986 230294
rect 552222 230058 552306 230294
rect 552542 230058 552574 230294
rect 551954 194614 552574 230058
rect 551954 194378 551986 194614
rect 552222 194378 552306 194614
rect 552542 194378 552574 194614
rect 551954 194294 552574 194378
rect 551954 194058 551986 194294
rect 552222 194058 552306 194294
rect 552542 194058 552574 194294
rect 551954 158614 552574 194058
rect 551954 158378 551986 158614
rect 552222 158378 552306 158614
rect 552542 158378 552574 158614
rect 551954 158294 552574 158378
rect 551954 158058 551986 158294
rect 552222 158058 552306 158294
rect 552542 158058 552574 158294
rect 551954 122614 552574 158058
rect 551954 122378 551986 122614
rect 552222 122378 552306 122614
rect 552542 122378 552574 122614
rect 551954 122294 552574 122378
rect 551954 122058 551986 122294
rect 552222 122058 552306 122294
rect 552542 122058 552574 122294
rect 551954 86614 552574 122058
rect 551954 86378 551986 86614
rect 552222 86378 552306 86614
rect 552542 86378 552574 86614
rect 551954 86294 552574 86378
rect 551954 86058 551986 86294
rect 552222 86058 552306 86294
rect 552542 86058 552574 86294
rect 551954 50614 552574 86058
rect 551954 50378 551986 50614
rect 552222 50378 552306 50614
rect 552542 50378 552574 50614
rect 551954 50294 552574 50378
rect 551954 50058 551986 50294
rect 552222 50058 552306 50294
rect 552542 50058 552574 50294
rect 551954 14614 552574 50058
rect 551954 14378 551986 14614
rect 552222 14378 552306 14614
rect 552542 14378 552574 14614
rect 551954 14294 552574 14378
rect 551954 14058 551986 14294
rect 552222 14058 552306 14294
rect 552542 14058 552574 14294
rect 548234 -4422 548266 -4186
rect 548502 -4422 548586 -4186
rect 548822 -4422 548854 -4186
rect 548234 -4506 548854 -4422
rect 548234 -4742 548266 -4506
rect 548502 -4742 548586 -4506
rect 548822 -4742 548854 -4506
rect 548234 -5734 548854 -4742
rect 541954 -7302 541986 -7066
rect 542222 -7302 542306 -7066
rect 542542 -7302 542574 -7066
rect 541954 -7386 542574 -7302
rect 541954 -7622 541986 -7386
rect 542222 -7622 542306 -7386
rect 542542 -7622 542574 -7386
rect 541954 -7654 542574 -7622
rect 551954 -6106 552574 14058
rect 554514 707718 555134 707750
rect 554514 707482 554546 707718
rect 554782 707482 554866 707718
rect 555102 707482 555134 707718
rect 554514 707398 555134 707482
rect 554514 707162 554546 707398
rect 554782 707162 554866 707398
rect 555102 707162 555134 707398
rect 554514 673174 555134 707162
rect 554514 672938 554546 673174
rect 554782 672938 554866 673174
rect 555102 672938 555134 673174
rect 554514 672854 555134 672938
rect 554514 672618 554546 672854
rect 554782 672618 554866 672854
rect 555102 672618 555134 672854
rect 554514 637174 555134 672618
rect 554514 636938 554546 637174
rect 554782 636938 554866 637174
rect 555102 636938 555134 637174
rect 554514 636854 555134 636938
rect 554514 636618 554546 636854
rect 554782 636618 554866 636854
rect 555102 636618 555134 636854
rect 554514 601174 555134 636618
rect 554514 600938 554546 601174
rect 554782 600938 554866 601174
rect 555102 600938 555134 601174
rect 554514 600854 555134 600938
rect 554514 600618 554546 600854
rect 554782 600618 554866 600854
rect 555102 600618 555134 600854
rect 554514 565174 555134 600618
rect 554514 564938 554546 565174
rect 554782 564938 554866 565174
rect 555102 564938 555134 565174
rect 554514 564854 555134 564938
rect 554514 564618 554546 564854
rect 554782 564618 554866 564854
rect 555102 564618 555134 564854
rect 554514 529174 555134 564618
rect 554514 528938 554546 529174
rect 554782 528938 554866 529174
rect 555102 528938 555134 529174
rect 554514 528854 555134 528938
rect 554514 528618 554546 528854
rect 554782 528618 554866 528854
rect 555102 528618 555134 528854
rect 554514 493174 555134 528618
rect 554514 492938 554546 493174
rect 554782 492938 554866 493174
rect 555102 492938 555134 493174
rect 554514 492854 555134 492938
rect 554514 492618 554546 492854
rect 554782 492618 554866 492854
rect 555102 492618 555134 492854
rect 554514 457174 555134 492618
rect 554514 456938 554546 457174
rect 554782 456938 554866 457174
rect 555102 456938 555134 457174
rect 554514 456854 555134 456938
rect 554514 456618 554546 456854
rect 554782 456618 554866 456854
rect 555102 456618 555134 456854
rect 554514 421174 555134 456618
rect 554514 420938 554546 421174
rect 554782 420938 554866 421174
rect 555102 420938 555134 421174
rect 554514 420854 555134 420938
rect 554514 420618 554546 420854
rect 554782 420618 554866 420854
rect 555102 420618 555134 420854
rect 554514 385174 555134 420618
rect 554514 384938 554546 385174
rect 554782 384938 554866 385174
rect 555102 384938 555134 385174
rect 554514 384854 555134 384938
rect 554514 384618 554546 384854
rect 554782 384618 554866 384854
rect 555102 384618 555134 384854
rect 554514 349174 555134 384618
rect 554514 348938 554546 349174
rect 554782 348938 554866 349174
rect 555102 348938 555134 349174
rect 554514 348854 555134 348938
rect 554514 348618 554546 348854
rect 554782 348618 554866 348854
rect 555102 348618 555134 348854
rect 554514 313174 555134 348618
rect 554514 312938 554546 313174
rect 554782 312938 554866 313174
rect 555102 312938 555134 313174
rect 554514 312854 555134 312938
rect 554514 312618 554546 312854
rect 554782 312618 554866 312854
rect 555102 312618 555134 312854
rect 554514 277174 555134 312618
rect 554514 276938 554546 277174
rect 554782 276938 554866 277174
rect 555102 276938 555134 277174
rect 554514 276854 555134 276938
rect 554514 276618 554546 276854
rect 554782 276618 554866 276854
rect 555102 276618 555134 276854
rect 554514 241174 555134 276618
rect 554514 240938 554546 241174
rect 554782 240938 554866 241174
rect 555102 240938 555134 241174
rect 554514 240854 555134 240938
rect 554514 240618 554546 240854
rect 554782 240618 554866 240854
rect 555102 240618 555134 240854
rect 554514 205174 555134 240618
rect 554514 204938 554546 205174
rect 554782 204938 554866 205174
rect 555102 204938 555134 205174
rect 554514 204854 555134 204938
rect 554514 204618 554546 204854
rect 554782 204618 554866 204854
rect 555102 204618 555134 204854
rect 554514 169174 555134 204618
rect 554514 168938 554546 169174
rect 554782 168938 554866 169174
rect 555102 168938 555134 169174
rect 554514 168854 555134 168938
rect 554514 168618 554546 168854
rect 554782 168618 554866 168854
rect 555102 168618 555134 168854
rect 554514 133174 555134 168618
rect 554514 132938 554546 133174
rect 554782 132938 554866 133174
rect 555102 132938 555134 133174
rect 554514 132854 555134 132938
rect 554514 132618 554546 132854
rect 554782 132618 554866 132854
rect 555102 132618 555134 132854
rect 554514 97174 555134 132618
rect 554514 96938 554546 97174
rect 554782 96938 554866 97174
rect 555102 96938 555134 97174
rect 554514 96854 555134 96938
rect 554514 96618 554546 96854
rect 554782 96618 554866 96854
rect 555102 96618 555134 96854
rect 554514 61174 555134 96618
rect 554514 60938 554546 61174
rect 554782 60938 554866 61174
rect 555102 60938 555134 61174
rect 554514 60854 555134 60938
rect 554514 60618 554546 60854
rect 554782 60618 554866 60854
rect 555102 60618 555134 60854
rect 554514 25174 555134 60618
rect 554514 24938 554546 25174
rect 554782 24938 554866 25174
rect 555102 24938 555134 25174
rect 554514 24854 555134 24938
rect 554514 24618 554546 24854
rect 554782 24618 554866 24854
rect 555102 24618 555134 24854
rect 554514 -3226 555134 24618
rect 554514 -3462 554546 -3226
rect 554782 -3462 554866 -3226
rect 555102 -3462 555134 -3226
rect 554514 -3546 555134 -3462
rect 554514 -3782 554546 -3546
rect 554782 -3782 554866 -3546
rect 555102 -3782 555134 -3546
rect 554514 -3814 555134 -3782
rect 558234 676894 558854 709082
rect 558234 676658 558266 676894
rect 558502 676658 558586 676894
rect 558822 676658 558854 676894
rect 558234 676574 558854 676658
rect 558234 676338 558266 676574
rect 558502 676338 558586 676574
rect 558822 676338 558854 676574
rect 558234 640894 558854 676338
rect 558234 640658 558266 640894
rect 558502 640658 558586 640894
rect 558822 640658 558854 640894
rect 558234 640574 558854 640658
rect 558234 640338 558266 640574
rect 558502 640338 558586 640574
rect 558822 640338 558854 640574
rect 558234 604894 558854 640338
rect 558234 604658 558266 604894
rect 558502 604658 558586 604894
rect 558822 604658 558854 604894
rect 558234 604574 558854 604658
rect 558234 604338 558266 604574
rect 558502 604338 558586 604574
rect 558822 604338 558854 604574
rect 558234 568894 558854 604338
rect 558234 568658 558266 568894
rect 558502 568658 558586 568894
rect 558822 568658 558854 568894
rect 558234 568574 558854 568658
rect 558234 568338 558266 568574
rect 558502 568338 558586 568574
rect 558822 568338 558854 568574
rect 558234 532894 558854 568338
rect 558234 532658 558266 532894
rect 558502 532658 558586 532894
rect 558822 532658 558854 532894
rect 558234 532574 558854 532658
rect 558234 532338 558266 532574
rect 558502 532338 558586 532574
rect 558822 532338 558854 532574
rect 558234 496894 558854 532338
rect 558234 496658 558266 496894
rect 558502 496658 558586 496894
rect 558822 496658 558854 496894
rect 558234 496574 558854 496658
rect 558234 496338 558266 496574
rect 558502 496338 558586 496574
rect 558822 496338 558854 496574
rect 558234 460894 558854 496338
rect 558234 460658 558266 460894
rect 558502 460658 558586 460894
rect 558822 460658 558854 460894
rect 558234 460574 558854 460658
rect 558234 460338 558266 460574
rect 558502 460338 558586 460574
rect 558822 460338 558854 460574
rect 558234 424894 558854 460338
rect 558234 424658 558266 424894
rect 558502 424658 558586 424894
rect 558822 424658 558854 424894
rect 558234 424574 558854 424658
rect 558234 424338 558266 424574
rect 558502 424338 558586 424574
rect 558822 424338 558854 424574
rect 558234 388894 558854 424338
rect 558234 388658 558266 388894
rect 558502 388658 558586 388894
rect 558822 388658 558854 388894
rect 558234 388574 558854 388658
rect 558234 388338 558266 388574
rect 558502 388338 558586 388574
rect 558822 388338 558854 388574
rect 558234 352894 558854 388338
rect 558234 352658 558266 352894
rect 558502 352658 558586 352894
rect 558822 352658 558854 352894
rect 558234 352574 558854 352658
rect 558234 352338 558266 352574
rect 558502 352338 558586 352574
rect 558822 352338 558854 352574
rect 558234 316894 558854 352338
rect 558234 316658 558266 316894
rect 558502 316658 558586 316894
rect 558822 316658 558854 316894
rect 558234 316574 558854 316658
rect 558234 316338 558266 316574
rect 558502 316338 558586 316574
rect 558822 316338 558854 316574
rect 558234 280894 558854 316338
rect 558234 280658 558266 280894
rect 558502 280658 558586 280894
rect 558822 280658 558854 280894
rect 558234 280574 558854 280658
rect 558234 280338 558266 280574
rect 558502 280338 558586 280574
rect 558822 280338 558854 280574
rect 558234 244894 558854 280338
rect 558234 244658 558266 244894
rect 558502 244658 558586 244894
rect 558822 244658 558854 244894
rect 558234 244574 558854 244658
rect 558234 244338 558266 244574
rect 558502 244338 558586 244574
rect 558822 244338 558854 244574
rect 558234 208894 558854 244338
rect 558234 208658 558266 208894
rect 558502 208658 558586 208894
rect 558822 208658 558854 208894
rect 558234 208574 558854 208658
rect 558234 208338 558266 208574
rect 558502 208338 558586 208574
rect 558822 208338 558854 208574
rect 558234 172894 558854 208338
rect 558234 172658 558266 172894
rect 558502 172658 558586 172894
rect 558822 172658 558854 172894
rect 558234 172574 558854 172658
rect 558234 172338 558266 172574
rect 558502 172338 558586 172574
rect 558822 172338 558854 172574
rect 558234 136894 558854 172338
rect 558234 136658 558266 136894
rect 558502 136658 558586 136894
rect 558822 136658 558854 136894
rect 558234 136574 558854 136658
rect 558234 136338 558266 136574
rect 558502 136338 558586 136574
rect 558822 136338 558854 136574
rect 558234 100894 558854 136338
rect 558234 100658 558266 100894
rect 558502 100658 558586 100894
rect 558822 100658 558854 100894
rect 558234 100574 558854 100658
rect 558234 100338 558266 100574
rect 558502 100338 558586 100574
rect 558822 100338 558854 100574
rect 558234 64894 558854 100338
rect 558234 64658 558266 64894
rect 558502 64658 558586 64894
rect 558822 64658 558854 64894
rect 558234 64574 558854 64658
rect 558234 64338 558266 64574
rect 558502 64338 558586 64574
rect 558822 64338 558854 64574
rect 558234 28894 558854 64338
rect 558234 28658 558266 28894
rect 558502 28658 558586 28894
rect 558822 28658 558854 28894
rect 558234 28574 558854 28658
rect 558234 28338 558266 28574
rect 558502 28338 558586 28574
rect 558822 28338 558854 28574
rect 558234 -5146 558854 28338
rect 560794 704838 561414 705830
rect 560794 704602 560826 704838
rect 561062 704602 561146 704838
rect 561382 704602 561414 704838
rect 560794 704518 561414 704602
rect 560794 704282 560826 704518
rect 561062 704282 561146 704518
rect 561382 704282 561414 704518
rect 560794 687454 561414 704282
rect 560794 687218 560826 687454
rect 561062 687218 561146 687454
rect 561382 687218 561414 687454
rect 560794 687134 561414 687218
rect 560794 686898 560826 687134
rect 561062 686898 561146 687134
rect 561382 686898 561414 687134
rect 560794 651454 561414 686898
rect 560794 651218 560826 651454
rect 561062 651218 561146 651454
rect 561382 651218 561414 651454
rect 560794 651134 561414 651218
rect 560794 650898 560826 651134
rect 561062 650898 561146 651134
rect 561382 650898 561414 651134
rect 560794 615454 561414 650898
rect 560794 615218 560826 615454
rect 561062 615218 561146 615454
rect 561382 615218 561414 615454
rect 560794 615134 561414 615218
rect 560794 614898 560826 615134
rect 561062 614898 561146 615134
rect 561382 614898 561414 615134
rect 560794 579454 561414 614898
rect 560794 579218 560826 579454
rect 561062 579218 561146 579454
rect 561382 579218 561414 579454
rect 560794 579134 561414 579218
rect 560794 578898 560826 579134
rect 561062 578898 561146 579134
rect 561382 578898 561414 579134
rect 560794 543454 561414 578898
rect 560794 543218 560826 543454
rect 561062 543218 561146 543454
rect 561382 543218 561414 543454
rect 560794 543134 561414 543218
rect 560794 542898 560826 543134
rect 561062 542898 561146 543134
rect 561382 542898 561414 543134
rect 560794 507454 561414 542898
rect 560794 507218 560826 507454
rect 561062 507218 561146 507454
rect 561382 507218 561414 507454
rect 560794 507134 561414 507218
rect 560794 506898 560826 507134
rect 561062 506898 561146 507134
rect 561382 506898 561414 507134
rect 560794 471454 561414 506898
rect 560794 471218 560826 471454
rect 561062 471218 561146 471454
rect 561382 471218 561414 471454
rect 560794 471134 561414 471218
rect 560794 470898 560826 471134
rect 561062 470898 561146 471134
rect 561382 470898 561414 471134
rect 560794 435454 561414 470898
rect 560794 435218 560826 435454
rect 561062 435218 561146 435454
rect 561382 435218 561414 435454
rect 560794 435134 561414 435218
rect 560794 434898 560826 435134
rect 561062 434898 561146 435134
rect 561382 434898 561414 435134
rect 560794 399454 561414 434898
rect 560794 399218 560826 399454
rect 561062 399218 561146 399454
rect 561382 399218 561414 399454
rect 560794 399134 561414 399218
rect 560794 398898 560826 399134
rect 561062 398898 561146 399134
rect 561382 398898 561414 399134
rect 560794 363454 561414 398898
rect 560794 363218 560826 363454
rect 561062 363218 561146 363454
rect 561382 363218 561414 363454
rect 560794 363134 561414 363218
rect 560794 362898 560826 363134
rect 561062 362898 561146 363134
rect 561382 362898 561414 363134
rect 560794 327454 561414 362898
rect 560794 327218 560826 327454
rect 561062 327218 561146 327454
rect 561382 327218 561414 327454
rect 560794 327134 561414 327218
rect 560794 326898 560826 327134
rect 561062 326898 561146 327134
rect 561382 326898 561414 327134
rect 560794 291454 561414 326898
rect 560794 291218 560826 291454
rect 561062 291218 561146 291454
rect 561382 291218 561414 291454
rect 560794 291134 561414 291218
rect 560794 290898 560826 291134
rect 561062 290898 561146 291134
rect 561382 290898 561414 291134
rect 560794 255454 561414 290898
rect 560794 255218 560826 255454
rect 561062 255218 561146 255454
rect 561382 255218 561414 255454
rect 560794 255134 561414 255218
rect 560794 254898 560826 255134
rect 561062 254898 561146 255134
rect 561382 254898 561414 255134
rect 560794 219454 561414 254898
rect 560794 219218 560826 219454
rect 561062 219218 561146 219454
rect 561382 219218 561414 219454
rect 560794 219134 561414 219218
rect 560794 218898 560826 219134
rect 561062 218898 561146 219134
rect 561382 218898 561414 219134
rect 560794 183454 561414 218898
rect 560794 183218 560826 183454
rect 561062 183218 561146 183454
rect 561382 183218 561414 183454
rect 560794 183134 561414 183218
rect 560794 182898 560826 183134
rect 561062 182898 561146 183134
rect 561382 182898 561414 183134
rect 560794 147454 561414 182898
rect 560794 147218 560826 147454
rect 561062 147218 561146 147454
rect 561382 147218 561414 147454
rect 560794 147134 561414 147218
rect 560794 146898 560826 147134
rect 561062 146898 561146 147134
rect 561382 146898 561414 147134
rect 560794 111454 561414 146898
rect 560794 111218 560826 111454
rect 561062 111218 561146 111454
rect 561382 111218 561414 111454
rect 560794 111134 561414 111218
rect 560794 110898 560826 111134
rect 561062 110898 561146 111134
rect 561382 110898 561414 111134
rect 560794 75454 561414 110898
rect 560794 75218 560826 75454
rect 561062 75218 561146 75454
rect 561382 75218 561414 75454
rect 560794 75134 561414 75218
rect 560794 74898 560826 75134
rect 561062 74898 561146 75134
rect 561382 74898 561414 75134
rect 560794 39454 561414 74898
rect 560794 39218 560826 39454
rect 561062 39218 561146 39454
rect 561382 39218 561414 39454
rect 560794 39134 561414 39218
rect 560794 38898 560826 39134
rect 561062 38898 561146 39134
rect 561382 38898 561414 39134
rect 560794 3454 561414 38898
rect 560794 3218 560826 3454
rect 561062 3218 561146 3454
rect 561382 3218 561414 3454
rect 560794 3134 561414 3218
rect 560794 2898 560826 3134
rect 561062 2898 561146 3134
rect 561382 2898 561414 3134
rect 560794 -346 561414 2898
rect 560794 -582 560826 -346
rect 561062 -582 561146 -346
rect 561382 -582 561414 -346
rect 560794 -666 561414 -582
rect 560794 -902 560826 -666
rect 561062 -902 561146 -666
rect 561382 -902 561414 -666
rect 560794 -1894 561414 -902
rect 561954 680614 562574 711002
rect 571954 710598 572574 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 571954 710362 571986 710598
rect 572222 710362 572306 710598
rect 572542 710362 572574 710598
rect 571954 710278 572574 710362
rect 571954 710042 571986 710278
rect 572222 710042 572306 710278
rect 572542 710042 572574 710278
rect 568234 708678 568854 709670
rect 568234 708442 568266 708678
rect 568502 708442 568586 708678
rect 568822 708442 568854 708678
rect 568234 708358 568854 708442
rect 568234 708122 568266 708358
rect 568502 708122 568586 708358
rect 568822 708122 568854 708358
rect 561954 680378 561986 680614
rect 562222 680378 562306 680614
rect 562542 680378 562574 680614
rect 561954 680294 562574 680378
rect 561954 680058 561986 680294
rect 562222 680058 562306 680294
rect 562542 680058 562574 680294
rect 561954 644614 562574 680058
rect 561954 644378 561986 644614
rect 562222 644378 562306 644614
rect 562542 644378 562574 644614
rect 561954 644294 562574 644378
rect 561954 644058 561986 644294
rect 562222 644058 562306 644294
rect 562542 644058 562574 644294
rect 561954 608614 562574 644058
rect 561954 608378 561986 608614
rect 562222 608378 562306 608614
rect 562542 608378 562574 608614
rect 561954 608294 562574 608378
rect 561954 608058 561986 608294
rect 562222 608058 562306 608294
rect 562542 608058 562574 608294
rect 561954 572614 562574 608058
rect 561954 572378 561986 572614
rect 562222 572378 562306 572614
rect 562542 572378 562574 572614
rect 561954 572294 562574 572378
rect 561954 572058 561986 572294
rect 562222 572058 562306 572294
rect 562542 572058 562574 572294
rect 561954 536614 562574 572058
rect 561954 536378 561986 536614
rect 562222 536378 562306 536614
rect 562542 536378 562574 536614
rect 561954 536294 562574 536378
rect 561954 536058 561986 536294
rect 562222 536058 562306 536294
rect 562542 536058 562574 536294
rect 561954 500614 562574 536058
rect 561954 500378 561986 500614
rect 562222 500378 562306 500614
rect 562542 500378 562574 500614
rect 561954 500294 562574 500378
rect 561954 500058 561986 500294
rect 562222 500058 562306 500294
rect 562542 500058 562574 500294
rect 561954 464614 562574 500058
rect 561954 464378 561986 464614
rect 562222 464378 562306 464614
rect 562542 464378 562574 464614
rect 561954 464294 562574 464378
rect 561954 464058 561986 464294
rect 562222 464058 562306 464294
rect 562542 464058 562574 464294
rect 561954 428614 562574 464058
rect 561954 428378 561986 428614
rect 562222 428378 562306 428614
rect 562542 428378 562574 428614
rect 561954 428294 562574 428378
rect 561954 428058 561986 428294
rect 562222 428058 562306 428294
rect 562542 428058 562574 428294
rect 561954 392614 562574 428058
rect 561954 392378 561986 392614
rect 562222 392378 562306 392614
rect 562542 392378 562574 392614
rect 561954 392294 562574 392378
rect 561954 392058 561986 392294
rect 562222 392058 562306 392294
rect 562542 392058 562574 392294
rect 561954 356614 562574 392058
rect 561954 356378 561986 356614
rect 562222 356378 562306 356614
rect 562542 356378 562574 356614
rect 561954 356294 562574 356378
rect 561954 356058 561986 356294
rect 562222 356058 562306 356294
rect 562542 356058 562574 356294
rect 561954 320614 562574 356058
rect 561954 320378 561986 320614
rect 562222 320378 562306 320614
rect 562542 320378 562574 320614
rect 561954 320294 562574 320378
rect 561954 320058 561986 320294
rect 562222 320058 562306 320294
rect 562542 320058 562574 320294
rect 561954 284614 562574 320058
rect 561954 284378 561986 284614
rect 562222 284378 562306 284614
rect 562542 284378 562574 284614
rect 561954 284294 562574 284378
rect 561954 284058 561986 284294
rect 562222 284058 562306 284294
rect 562542 284058 562574 284294
rect 561954 248614 562574 284058
rect 561954 248378 561986 248614
rect 562222 248378 562306 248614
rect 562542 248378 562574 248614
rect 561954 248294 562574 248378
rect 561954 248058 561986 248294
rect 562222 248058 562306 248294
rect 562542 248058 562574 248294
rect 561954 212614 562574 248058
rect 561954 212378 561986 212614
rect 562222 212378 562306 212614
rect 562542 212378 562574 212614
rect 561954 212294 562574 212378
rect 561954 212058 561986 212294
rect 562222 212058 562306 212294
rect 562542 212058 562574 212294
rect 561954 176614 562574 212058
rect 561954 176378 561986 176614
rect 562222 176378 562306 176614
rect 562542 176378 562574 176614
rect 561954 176294 562574 176378
rect 561954 176058 561986 176294
rect 562222 176058 562306 176294
rect 562542 176058 562574 176294
rect 561954 140614 562574 176058
rect 561954 140378 561986 140614
rect 562222 140378 562306 140614
rect 562542 140378 562574 140614
rect 561954 140294 562574 140378
rect 561954 140058 561986 140294
rect 562222 140058 562306 140294
rect 562542 140058 562574 140294
rect 561954 104614 562574 140058
rect 561954 104378 561986 104614
rect 562222 104378 562306 104614
rect 562542 104378 562574 104614
rect 561954 104294 562574 104378
rect 561954 104058 561986 104294
rect 562222 104058 562306 104294
rect 562542 104058 562574 104294
rect 561954 68614 562574 104058
rect 561954 68378 561986 68614
rect 562222 68378 562306 68614
rect 562542 68378 562574 68614
rect 561954 68294 562574 68378
rect 561954 68058 561986 68294
rect 562222 68058 562306 68294
rect 562542 68058 562574 68294
rect 561954 32614 562574 68058
rect 561954 32378 561986 32614
rect 562222 32378 562306 32614
rect 562542 32378 562574 32614
rect 561954 32294 562574 32378
rect 561954 32058 561986 32294
rect 562222 32058 562306 32294
rect 562542 32058 562574 32294
rect 558234 -5382 558266 -5146
rect 558502 -5382 558586 -5146
rect 558822 -5382 558854 -5146
rect 558234 -5466 558854 -5382
rect 558234 -5702 558266 -5466
rect 558502 -5702 558586 -5466
rect 558822 -5702 558854 -5466
rect 558234 -5734 558854 -5702
rect 551954 -6342 551986 -6106
rect 552222 -6342 552306 -6106
rect 552542 -6342 552574 -6106
rect 551954 -6426 552574 -6342
rect 551954 -6662 551986 -6426
rect 552222 -6662 552306 -6426
rect 552542 -6662 552574 -6426
rect 551954 -7654 552574 -6662
rect 561954 -7066 562574 32058
rect 564514 706758 565134 707750
rect 564514 706522 564546 706758
rect 564782 706522 564866 706758
rect 565102 706522 565134 706758
rect 564514 706438 565134 706522
rect 564514 706202 564546 706438
rect 564782 706202 564866 706438
rect 565102 706202 565134 706438
rect 564514 691174 565134 706202
rect 564514 690938 564546 691174
rect 564782 690938 564866 691174
rect 565102 690938 565134 691174
rect 564514 690854 565134 690938
rect 564514 690618 564546 690854
rect 564782 690618 564866 690854
rect 565102 690618 565134 690854
rect 564514 655174 565134 690618
rect 564514 654938 564546 655174
rect 564782 654938 564866 655174
rect 565102 654938 565134 655174
rect 564514 654854 565134 654938
rect 564514 654618 564546 654854
rect 564782 654618 564866 654854
rect 565102 654618 565134 654854
rect 564514 619174 565134 654618
rect 564514 618938 564546 619174
rect 564782 618938 564866 619174
rect 565102 618938 565134 619174
rect 564514 618854 565134 618938
rect 564514 618618 564546 618854
rect 564782 618618 564866 618854
rect 565102 618618 565134 618854
rect 564514 583174 565134 618618
rect 564514 582938 564546 583174
rect 564782 582938 564866 583174
rect 565102 582938 565134 583174
rect 564514 582854 565134 582938
rect 564514 582618 564546 582854
rect 564782 582618 564866 582854
rect 565102 582618 565134 582854
rect 564514 547174 565134 582618
rect 564514 546938 564546 547174
rect 564782 546938 564866 547174
rect 565102 546938 565134 547174
rect 564514 546854 565134 546938
rect 564514 546618 564546 546854
rect 564782 546618 564866 546854
rect 565102 546618 565134 546854
rect 564514 511174 565134 546618
rect 564514 510938 564546 511174
rect 564782 510938 564866 511174
rect 565102 510938 565134 511174
rect 564514 510854 565134 510938
rect 564514 510618 564546 510854
rect 564782 510618 564866 510854
rect 565102 510618 565134 510854
rect 564514 475174 565134 510618
rect 564514 474938 564546 475174
rect 564782 474938 564866 475174
rect 565102 474938 565134 475174
rect 564514 474854 565134 474938
rect 564514 474618 564546 474854
rect 564782 474618 564866 474854
rect 565102 474618 565134 474854
rect 564514 439174 565134 474618
rect 564514 438938 564546 439174
rect 564782 438938 564866 439174
rect 565102 438938 565134 439174
rect 564514 438854 565134 438938
rect 564514 438618 564546 438854
rect 564782 438618 564866 438854
rect 565102 438618 565134 438854
rect 564514 403174 565134 438618
rect 564514 402938 564546 403174
rect 564782 402938 564866 403174
rect 565102 402938 565134 403174
rect 564514 402854 565134 402938
rect 564514 402618 564546 402854
rect 564782 402618 564866 402854
rect 565102 402618 565134 402854
rect 564514 367174 565134 402618
rect 564514 366938 564546 367174
rect 564782 366938 564866 367174
rect 565102 366938 565134 367174
rect 564514 366854 565134 366938
rect 564514 366618 564546 366854
rect 564782 366618 564866 366854
rect 565102 366618 565134 366854
rect 564514 331174 565134 366618
rect 564514 330938 564546 331174
rect 564782 330938 564866 331174
rect 565102 330938 565134 331174
rect 564514 330854 565134 330938
rect 564514 330618 564546 330854
rect 564782 330618 564866 330854
rect 565102 330618 565134 330854
rect 564514 295174 565134 330618
rect 564514 294938 564546 295174
rect 564782 294938 564866 295174
rect 565102 294938 565134 295174
rect 564514 294854 565134 294938
rect 564514 294618 564546 294854
rect 564782 294618 564866 294854
rect 565102 294618 565134 294854
rect 564514 259174 565134 294618
rect 564514 258938 564546 259174
rect 564782 258938 564866 259174
rect 565102 258938 565134 259174
rect 564514 258854 565134 258938
rect 564514 258618 564546 258854
rect 564782 258618 564866 258854
rect 565102 258618 565134 258854
rect 564514 223174 565134 258618
rect 564514 222938 564546 223174
rect 564782 222938 564866 223174
rect 565102 222938 565134 223174
rect 564514 222854 565134 222938
rect 564514 222618 564546 222854
rect 564782 222618 564866 222854
rect 565102 222618 565134 222854
rect 564514 187174 565134 222618
rect 564514 186938 564546 187174
rect 564782 186938 564866 187174
rect 565102 186938 565134 187174
rect 564514 186854 565134 186938
rect 564514 186618 564546 186854
rect 564782 186618 564866 186854
rect 565102 186618 565134 186854
rect 564514 151174 565134 186618
rect 564514 150938 564546 151174
rect 564782 150938 564866 151174
rect 565102 150938 565134 151174
rect 564514 150854 565134 150938
rect 564514 150618 564546 150854
rect 564782 150618 564866 150854
rect 565102 150618 565134 150854
rect 564514 115174 565134 150618
rect 564514 114938 564546 115174
rect 564782 114938 564866 115174
rect 565102 114938 565134 115174
rect 564514 114854 565134 114938
rect 564514 114618 564546 114854
rect 564782 114618 564866 114854
rect 565102 114618 565134 114854
rect 564514 79174 565134 114618
rect 564514 78938 564546 79174
rect 564782 78938 564866 79174
rect 565102 78938 565134 79174
rect 564514 78854 565134 78938
rect 564514 78618 564546 78854
rect 564782 78618 564866 78854
rect 565102 78618 565134 78854
rect 564514 43174 565134 78618
rect 564514 42938 564546 43174
rect 564782 42938 564866 43174
rect 565102 42938 565134 43174
rect 564514 42854 565134 42938
rect 564514 42618 564546 42854
rect 564782 42618 564866 42854
rect 565102 42618 565134 42854
rect 564514 7174 565134 42618
rect 564514 6938 564546 7174
rect 564782 6938 564866 7174
rect 565102 6938 565134 7174
rect 564514 6854 565134 6938
rect 564514 6618 564546 6854
rect 564782 6618 564866 6854
rect 565102 6618 565134 6854
rect 564514 -2266 565134 6618
rect 564514 -2502 564546 -2266
rect 564782 -2502 564866 -2266
rect 565102 -2502 565134 -2266
rect 564514 -2586 565134 -2502
rect 564514 -2822 564546 -2586
rect 564782 -2822 564866 -2586
rect 565102 -2822 565134 -2586
rect 564514 -3814 565134 -2822
rect 568234 694894 568854 708122
rect 568234 694658 568266 694894
rect 568502 694658 568586 694894
rect 568822 694658 568854 694894
rect 568234 694574 568854 694658
rect 568234 694338 568266 694574
rect 568502 694338 568586 694574
rect 568822 694338 568854 694574
rect 568234 658894 568854 694338
rect 568234 658658 568266 658894
rect 568502 658658 568586 658894
rect 568822 658658 568854 658894
rect 568234 658574 568854 658658
rect 568234 658338 568266 658574
rect 568502 658338 568586 658574
rect 568822 658338 568854 658574
rect 568234 622894 568854 658338
rect 568234 622658 568266 622894
rect 568502 622658 568586 622894
rect 568822 622658 568854 622894
rect 568234 622574 568854 622658
rect 568234 622338 568266 622574
rect 568502 622338 568586 622574
rect 568822 622338 568854 622574
rect 568234 586894 568854 622338
rect 568234 586658 568266 586894
rect 568502 586658 568586 586894
rect 568822 586658 568854 586894
rect 568234 586574 568854 586658
rect 568234 586338 568266 586574
rect 568502 586338 568586 586574
rect 568822 586338 568854 586574
rect 568234 550894 568854 586338
rect 568234 550658 568266 550894
rect 568502 550658 568586 550894
rect 568822 550658 568854 550894
rect 568234 550574 568854 550658
rect 568234 550338 568266 550574
rect 568502 550338 568586 550574
rect 568822 550338 568854 550574
rect 568234 514894 568854 550338
rect 568234 514658 568266 514894
rect 568502 514658 568586 514894
rect 568822 514658 568854 514894
rect 568234 514574 568854 514658
rect 568234 514338 568266 514574
rect 568502 514338 568586 514574
rect 568822 514338 568854 514574
rect 568234 478894 568854 514338
rect 568234 478658 568266 478894
rect 568502 478658 568586 478894
rect 568822 478658 568854 478894
rect 568234 478574 568854 478658
rect 568234 478338 568266 478574
rect 568502 478338 568586 478574
rect 568822 478338 568854 478574
rect 568234 442894 568854 478338
rect 568234 442658 568266 442894
rect 568502 442658 568586 442894
rect 568822 442658 568854 442894
rect 568234 442574 568854 442658
rect 568234 442338 568266 442574
rect 568502 442338 568586 442574
rect 568822 442338 568854 442574
rect 568234 406894 568854 442338
rect 568234 406658 568266 406894
rect 568502 406658 568586 406894
rect 568822 406658 568854 406894
rect 568234 406574 568854 406658
rect 568234 406338 568266 406574
rect 568502 406338 568586 406574
rect 568822 406338 568854 406574
rect 568234 370894 568854 406338
rect 568234 370658 568266 370894
rect 568502 370658 568586 370894
rect 568822 370658 568854 370894
rect 568234 370574 568854 370658
rect 568234 370338 568266 370574
rect 568502 370338 568586 370574
rect 568822 370338 568854 370574
rect 568234 334894 568854 370338
rect 568234 334658 568266 334894
rect 568502 334658 568586 334894
rect 568822 334658 568854 334894
rect 568234 334574 568854 334658
rect 568234 334338 568266 334574
rect 568502 334338 568586 334574
rect 568822 334338 568854 334574
rect 568234 298894 568854 334338
rect 568234 298658 568266 298894
rect 568502 298658 568586 298894
rect 568822 298658 568854 298894
rect 568234 298574 568854 298658
rect 568234 298338 568266 298574
rect 568502 298338 568586 298574
rect 568822 298338 568854 298574
rect 568234 262894 568854 298338
rect 568234 262658 568266 262894
rect 568502 262658 568586 262894
rect 568822 262658 568854 262894
rect 568234 262574 568854 262658
rect 568234 262338 568266 262574
rect 568502 262338 568586 262574
rect 568822 262338 568854 262574
rect 568234 226894 568854 262338
rect 568234 226658 568266 226894
rect 568502 226658 568586 226894
rect 568822 226658 568854 226894
rect 568234 226574 568854 226658
rect 568234 226338 568266 226574
rect 568502 226338 568586 226574
rect 568822 226338 568854 226574
rect 568234 190894 568854 226338
rect 568234 190658 568266 190894
rect 568502 190658 568586 190894
rect 568822 190658 568854 190894
rect 568234 190574 568854 190658
rect 568234 190338 568266 190574
rect 568502 190338 568586 190574
rect 568822 190338 568854 190574
rect 568234 154894 568854 190338
rect 568234 154658 568266 154894
rect 568502 154658 568586 154894
rect 568822 154658 568854 154894
rect 568234 154574 568854 154658
rect 568234 154338 568266 154574
rect 568502 154338 568586 154574
rect 568822 154338 568854 154574
rect 568234 118894 568854 154338
rect 568234 118658 568266 118894
rect 568502 118658 568586 118894
rect 568822 118658 568854 118894
rect 568234 118574 568854 118658
rect 568234 118338 568266 118574
rect 568502 118338 568586 118574
rect 568822 118338 568854 118574
rect 568234 82894 568854 118338
rect 568234 82658 568266 82894
rect 568502 82658 568586 82894
rect 568822 82658 568854 82894
rect 568234 82574 568854 82658
rect 568234 82338 568266 82574
rect 568502 82338 568586 82574
rect 568822 82338 568854 82574
rect 568234 46894 568854 82338
rect 568234 46658 568266 46894
rect 568502 46658 568586 46894
rect 568822 46658 568854 46894
rect 568234 46574 568854 46658
rect 568234 46338 568266 46574
rect 568502 46338 568586 46574
rect 568822 46338 568854 46574
rect 568234 10894 568854 46338
rect 568234 10658 568266 10894
rect 568502 10658 568586 10894
rect 568822 10658 568854 10894
rect 568234 10574 568854 10658
rect 568234 10338 568266 10574
rect 568502 10338 568586 10574
rect 568822 10338 568854 10574
rect 568234 -4186 568854 10338
rect 570794 705798 571414 705830
rect 570794 705562 570826 705798
rect 571062 705562 571146 705798
rect 571382 705562 571414 705798
rect 570794 705478 571414 705562
rect 570794 705242 570826 705478
rect 571062 705242 571146 705478
rect 571382 705242 571414 705478
rect 570794 669454 571414 705242
rect 570794 669218 570826 669454
rect 571062 669218 571146 669454
rect 571382 669218 571414 669454
rect 570794 669134 571414 669218
rect 570794 668898 570826 669134
rect 571062 668898 571146 669134
rect 571382 668898 571414 669134
rect 570794 633454 571414 668898
rect 570794 633218 570826 633454
rect 571062 633218 571146 633454
rect 571382 633218 571414 633454
rect 570794 633134 571414 633218
rect 570794 632898 570826 633134
rect 571062 632898 571146 633134
rect 571382 632898 571414 633134
rect 570794 597454 571414 632898
rect 570794 597218 570826 597454
rect 571062 597218 571146 597454
rect 571382 597218 571414 597454
rect 570794 597134 571414 597218
rect 570794 596898 570826 597134
rect 571062 596898 571146 597134
rect 571382 596898 571414 597134
rect 570794 561454 571414 596898
rect 570794 561218 570826 561454
rect 571062 561218 571146 561454
rect 571382 561218 571414 561454
rect 570794 561134 571414 561218
rect 570794 560898 570826 561134
rect 571062 560898 571146 561134
rect 571382 560898 571414 561134
rect 570794 525454 571414 560898
rect 570794 525218 570826 525454
rect 571062 525218 571146 525454
rect 571382 525218 571414 525454
rect 570794 525134 571414 525218
rect 570794 524898 570826 525134
rect 571062 524898 571146 525134
rect 571382 524898 571414 525134
rect 570794 489454 571414 524898
rect 570794 489218 570826 489454
rect 571062 489218 571146 489454
rect 571382 489218 571414 489454
rect 570794 489134 571414 489218
rect 570794 488898 570826 489134
rect 571062 488898 571146 489134
rect 571382 488898 571414 489134
rect 570794 453454 571414 488898
rect 570794 453218 570826 453454
rect 571062 453218 571146 453454
rect 571382 453218 571414 453454
rect 570794 453134 571414 453218
rect 570794 452898 570826 453134
rect 571062 452898 571146 453134
rect 571382 452898 571414 453134
rect 570794 417454 571414 452898
rect 570794 417218 570826 417454
rect 571062 417218 571146 417454
rect 571382 417218 571414 417454
rect 570794 417134 571414 417218
rect 570794 416898 570826 417134
rect 571062 416898 571146 417134
rect 571382 416898 571414 417134
rect 570794 381454 571414 416898
rect 570794 381218 570826 381454
rect 571062 381218 571146 381454
rect 571382 381218 571414 381454
rect 570794 381134 571414 381218
rect 570794 380898 570826 381134
rect 571062 380898 571146 381134
rect 571382 380898 571414 381134
rect 570794 345454 571414 380898
rect 570794 345218 570826 345454
rect 571062 345218 571146 345454
rect 571382 345218 571414 345454
rect 570794 345134 571414 345218
rect 570794 344898 570826 345134
rect 571062 344898 571146 345134
rect 571382 344898 571414 345134
rect 570794 309454 571414 344898
rect 570794 309218 570826 309454
rect 571062 309218 571146 309454
rect 571382 309218 571414 309454
rect 570794 309134 571414 309218
rect 570794 308898 570826 309134
rect 571062 308898 571146 309134
rect 571382 308898 571414 309134
rect 570794 273454 571414 308898
rect 570794 273218 570826 273454
rect 571062 273218 571146 273454
rect 571382 273218 571414 273454
rect 570794 273134 571414 273218
rect 570794 272898 570826 273134
rect 571062 272898 571146 273134
rect 571382 272898 571414 273134
rect 570794 237454 571414 272898
rect 570794 237218 570826 237454
rect 571062 237218 571146 237454
rect 571382 237218 571414 237454
rect 570794 237134 571414 237218
rect 570794 236898 570826 237134
rect 571062 236898 571146 237134
rect 571382 236898 571414 237134
rect 570794 201454 571414 236898
rect 570794 201218 570826 201454
rect 571062 201218 571146 201454
rect 571382 201218 571414 201454
rect 570794 201134 571414 201218
rect 570794 200898 570826 201134
rect 571062 200898 571146 201134
rect 571382 200898 571414 201134
rect 570794 165454 571414 200898
rect 570794 165218 570826 165454
rect 571062 165218 571146 165454
rect 571382 165218 571414 165454
rect 570794 165134 571414 165218
rect 570794 164898 570826 165134
rect 571062 164898 571146 165134
rect 571382 164898 571414 165134
rect 570794 129454 571414 164898
rect 570794 129218 570826 129454
rect 571062 129218 571146 129454
rect 571382 129218 571414 129454
rect 570794 129134 571414 129218
rect 570794 128898 570826 129134
rect 571062 128898 571146 129134
rect 571382 128898 571414 129134
rect 570794 93454 571414 128898
rect 570794 93218 570826 93454
rect 571062 93218 571146 93454
rect 571382 93218 571414 93454
rect 570794 93134 571414 93218
rect 570794 92898 570826 93134
rect 571062 92898 571146 93134
rect 571382 92898 571414 93134
rect 570794 57454 571414 92898
rect 570794 57218 570826 57454
rect 571062 57218 571146 57454
rect 571382 57218 571414 57454
rect 570794 57134 571414 57218
rect 570794 56898 570826 57134
rect 571062 56898 571146 57134
rect 571382 56898 571414 57134
rect 570794 21454 571414 56898
rect 570794 21218 570826 21454
rect 571062 21218 571146 21454
rect 571382 21218 571414 21454
rect 570794 21134 571414 21218
rect 570794 20898 570826 21134
rect 571062 20898 571146 21134
rect 571382 20898 571414 21134
rect 570794 -1306 571414 20898
rect 570794 -1542 570826 -1306
rect 571062 -1542 571146 -1306
rect 571382 -1542 571414 -1306
rect 570794 -1626 571414 -1542
rect 570794 -1862 570826 -1626
rect 571062 -1862 571146 -1626
rect 571382 -1862 571414 -1626
rect 570794 -1894 571414 -1862
rect 571954 698614 572574 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 578234 709638 578854 709670
rect 578234 709402 578266 709638
rect 578502 709402 578586 709638
rect 578822 709402 578854 709638
rect 578234 709318 578854 709402
rect 578234 709082 578266 709318
rect 578502 709082 578586 709318
rect 578822 709082 578854 709318
rect 571954 698378 571986 698614
rect 572222 698378 572306 698614
rect 572542 698378 572574 698614
rect 571954 698294 572574 698378
rect 571954 698058 571986 698294
rect 572222 698058 572306 698294
rect 572542 698058 572574 698294
rect 571954 662614 572574 698058
rect 571954 662378 571986 662614
rect 572222 662378 572306 662614
rect 572542 662378 572574 662614
rect 571954 662294 572574 662378
rect 571954 662058 571986 662294
rect 572222 662058 572306 662294
rect 572542 662058 572574 662294
rect 571954 626614 572574 662058
rect 571954 626378 571986 626614
rect 572222 626378 572306 626614
rect 572542 626378 572574 626614
rect 571954 626294 572574 626378
rect 571954 626058 571986 626294
rect 572222 626058 572306 626294
rect 572542 626058 572574 626294
rect 571954 590614 572574 626058
rect 571954 590378 571986 590614
rect 572222 590378 572306 590614
rect 572542 590378 572574 590614
rect 571954 590294 572574 590378
rect 571954 590058 571986 590294
rect 572222 590058 572306 590294
rect 572542 590058 572574 590294
rect 571954 554614 572574 590058
rect 571954 554378 571986 554614
rect 572222 554378 572306 554614
rect 572542 554378 572574 554614
rect 571954 554294 572574 554378
rect 571954 554058 571986 554294
rect 572222 554058 572306 554294
rect 572542 554058 572574 554294
rect 571954 518614 572574 554058
rect 571954 518378 571986 518614
rect 572222 518378 572306 518614
rect 572542 518378 572574 518614
rect 571954 518294 572574 518378
rect 571954 518058 571986 518294
rect 572222 518058 572306 518294
rect 572542 518058 572574 518294
rect 571954 482614 572574 518058
rect 571954 482378 571986 482614
rect 572222 482378 572306 482614
rect 572542 482378 572574 482614
rect 571954 482294 572574 482378
rect 571954 482058 571986 482294
rect 572222 482058 572306 482294
rect 572542 482058 572574 482294
rect 571954 446614 572574 482058
rect 571954 446378 571986 446614
rect 572222 446378 572306 446614
rect 572542 446378 572574 446614
rect 571954 446294 572574 446378
rect 571954 446058 571986 446294
rect 572222 446058 572306 446294
rect 572542 446058 572574 446294
rect 571954 410614 572574 446058
rect 571954 410378 571986 410614
rect 572222 410378 572306 410614
rect 572542 410378 572574 410614
rect 571954 410294 572574 410378
rect 571954 410058 571986 410294
rect 572222 410058 572306 410294
rect 572542 410058 572574 410294
rect 571954 374614 572574 410058
rect 571954 374378 571986 374614
rect 572222 374378 572306 374614
rect 572542 374378 572574 374614
rect 571954 374294 572574 374378
rect 571954 374058 571986 374294
rect 572222 374058 572306 374294
rect 572542 374058 572574 374294
rect 571954 338614 572574 374058
rect 571954 338378 571986 338614
rect 572222 338378 572306 338614
rect 572542 338378 572574 338614
rect 571954 338294 572574 338378
rect 571954 338058 571986 338294
rect 572222 338058 572306 338294
rect 572542 338058 572574 338294
rect 571954 302614 572574 338058
rect 571954 302378 571986 302614
rect 572222 302378 572306 302614
rect 572542 302378 572574 302614
rect 571954 302294 572574 302378
rect 571954 302058 571986 302294
rect 572222 302058 572306 302294
rect 572542 302058 572574 302294
rect 571954 266614 572574 302058
rect 571954 266378 571986 266614
rect 572222 266378 572306 266614
rect 572542 266378 572574 266614
rect 571954 266294 572574 266378
rect 571954 266058 571986 266294
rect 572222 266058 572306 266294
rect 572542 266058 572574 266294
rect 571954 230614 572574 266058
rect 571954 230378 571986 230614
rect 572222 230378 572306 230614
rect 572542 230378 572574 230614
rect 571954 230294 572574 230378
rect 571954 230058 571986 230294
rect 572222 230058 572306 230294
rect 572542 230058 572574 230294
rect 571954 194614 572574 230058
rect 571954 194378 571986 194614
rect 572222 194378 572306 194614
rect 572542 194378 572574 194614
rect 571954 194294 572574 194378
rect 571954 194058 571986 194294
rect 572222 194058 572306 194294
rect 572542 194058 572574 194294
rect 571954 158614 572574 194058
rect 571954 158378 571986 158614
rect 572222 158378 572306 158614
rect 572542 158378 572574 158614
rect 571954 158294 572574 158378
rect 571954 158058 571986 158294
rect 572222 158058 572306 158294
rect 572542 158058 572574 158294
rect 571954 122614 572574 158058
rect 571954 122378 571986 122614
rect 572222 122378 572306 122614
rect 572542 122378 572574 122614
rect 571954 122294 572574 122378
rect 571954 122058 571986 122294
rect 572222 122058 572306 122294
rect 572542 122058 572574 122294
rect 571954 86614 572574 122058
rect 571954 86378 571986 86614
rect 572222 86378 572306 86614
rect 572542 86378 572574 86614
rect 571954 86294 572574 86378
rect 571954 86058 571986 86294
rect 572222 86058 572306 86294
rect 572542 86058 572574 86294
rect 571954 50614 572574 86058
rect 571954 50378 571986 50614
rect 572222 50378 572306 50614
rect 572542 50378 572574 50614
rect 571954 50294 572574 50378
rect 571954 50058 571986 50294
rect 572222 50058 572306 50294
rect 572542 50058 572574 50294
rect 571954 14614 572574 50058
rect 571954 14378 571986 14614
rect 572222 14378 572306 14614
rect 572542 14378 572574 14614
rect 571954 14294 572574 14378
rect 571954 14058 571986 14294
rect 572222 14058 572306 14294
rect 572542 14058 572574 14294
rect 568234 -4422 568266 -4186
rect 568502 -4422 568586 -4186
rect 568822 -4422 568854 -4186
rect 568234 -4506 568854 -4422
rect 568234 -4742 568266 -4506
rect 568502 -4742 568586 -4506
rect 568822 -4742 568854 -4506
rect 568234 -5734 568854 -4742
rect 561954 -7302 561986 -7066
rect 562222 -7302 562306 -7066
rect 562542 -7302 562574 -7066
rect 561954 -7386 562574 -7302
rect 561954 -7622 561986 -7386
rect 562222 -7622 562306 -7386
rect 562542 -7622 562574 -7386
rect 561954 -7654 562574 -7622
rect 571954 -6106 572574 14058
rect 574514 707718 575134 707750
rect 574514 707482 574546 707718
rect 574782 707482 574866 707718
rect 575102 707482 575134 707718
rect 574514 707398 575134 707482
rect 574514 707162 574546 707398
rect 574782 707162 574866 707398
rect 575102 707162 575134 707398
rect 574514 673174 575134 707162
rect 574514 672938 574546 673174
rect 574782 672938 574866 673174
rect 575102 672938 575134 673174
rect 574514 672854 575134 672938
rect 574514 672618 574546 672854
rect 574782 672618 574866 672854
rect 575102 672618 575134 672854
rect 574514 637174 575134 672618
rect 574514 636938 574546 637174
rect 574782 636938 574866 637174
rect 575102 636938 575134 637174
rect 574514 636854 575134 636938
rect 574514 636618 574546 636854
rect 574782 636618 574866 636854
rect 575102 636618 575134 636854
rect 574514 601174 575134 636618
rect 574514 600938 574546 601174
rect 574782 600938 574866 601174
rect 575102 600938 575134 601174
rect 574514 600854 575134 600938
rect 574514 600618 574546 600854
rect 574782 600618 574866 600854
rect 575102 600618 575134 600854
rect 574514 565174 575134 600618
rect 574514 564938 574546 565174
rect 574782 564938 574866 565174
rect 575102 564938 575134 565174
rect 574514 564854 575134 564938
rect 574514 564618 574546 564854
rect 574782 564618 574866 564854
rect 575102 564618 575134 564854
rect 574514 529174 575134 564618
rect 574514 528938 574546 529174
rect 574782 528938 574866 529174
rect 575102 528938 575134 529174
rect 574514 528854 575134 528938
rect 574514 528618 574546 528854
rect 574782 528618 574866 528854
rect 575102 528618 575134 528854
rect 574514 493174 575134 528618
rect 574514 492938 574546 493174
rect 574782 492938 574866 493174
rect 575102 492938 575134 493174
rect 574514 492854 575134 492938
rect 574514 492618 574546 492854
rect 574782 492618 574866 492854
rect 575102 492618 575134 492854
rect 574514 457174 575134 492618
rect 574514 456938 574546 457174
rect 574782 456938 574866 457174
rect 575102 456938 575134 457174
rect 574514 456854 575134 456938
rect 574514 456618 574546 456854
rect 574782 456618 574866 456854
rect 575102 456618 575134 456854
rect 574514 421174 575134 456618
rect 574514 420938 574546 421174
rect 574782 420938 574866 421174
rect 575102 420938 575134 421174
rect 574514 420854 575134 420938
rect 574514 420618 574546 420854
rect 574782 420618 574866 420854
rect 575102 420618 575134 420854
rect 574514 385174 575134 420618
rect 574514 384938 574546 385174
rect 574782 384938 574866 385174
rect 575102 384938 575134 385174
rect 574514 384854 575134 384938
rect 574514 384618 574546 384854
rect 574782 384618 574866 384854
rect 575102 384618 575134 384854
rect 574514 349174 575134 384618
rect 574514 348938 574546 349174
rect 574782 348938 574866 349174
rect 575102 348938 575134 349174
rect 574514 348854 575134 348938
rect 574514 348618 574546 348854
rect 574782 348618 574866 348854
rect 575102 348618 575134 348854
rect 574514 313174 575134 348618
rect 574514 312938 574546 313174
rect 574782 312938 574866 313174
rect 575102 312938 575134 313174
rect 574514 312854 575134 312938
rect 574514 312618 574546 312854
rect 574782 312618 574866 312854
rect 575102 312618 575134 312854
rect 574514 277174 575134 312618
rect 574514 276938 574546 277174
rect 574782 276938 574866 277174
rect 575102 276938 575134 277174
rect 574514 276854 575134 276938
rect 574514 276618 574546 276854
rect 574782 276618 574866 276854
rect 575102 276618 575134 276854
rect 574514 241174 575134 276618
rect 574514 240938 574546 241174
rect 574782 240938 574866 241174
rect 575102 240938 575134 241174
rect 574514 240854 575134 240938
rect 574514 240618 574546 240854
rect 574782 240618 574866 240854
rect 575102 240618 575134 240854
rect 574514 205174 575134 240618
rect 574514 204938 574546 205174
rect 574782 204938 574866 205174
rect 575102 204938 575134 205174
rect 574514 204854 575134 204938
rect 574514 204618 574546 204854
rect 574782 204618 574866 204854
rect 575102 204618 575134 204854
rect 574514 169174 575134 204618
rect 574514 168938 574546 169174
rect 574782 168938 574866 169174
rect 575102 168938 575134 169174
rect 574514 168854 575134 168938
rect 574514 168618 574546 168854
rect 574782 168618 574866 168854
rect 575102 168618 575134 168854
rect 574514 133174 575134 168618
rect 574514 132938 574546 133174
rect 574782 132938 574866 133174
rect 575102 132938 575134 133174
rect 574514 132854 575134 132938
rect 574514 132618 574546 132854
rect 574782 132618 574866 132854
rect 575102 132618 575134 132854
rect 574514 97174 575134 132618
rect 574514 96938 574546 97174
rect 574782 96938 574866 97174
rect 575102 96938 575134 97174
rect 574514 96854 575134 96938
rect 574514 96618 574546 96854
rect 574782 96618 574866 96854
rect 575102 96618 575134 96854
rect 574514 61174 575134 96618
rect 574514 60938 574546 61174
rect 574782 60938 574866 61174
rect 575102 60938 575134 61174
rect 574514 60854 575134 60938
rect 574514 60618 574546 60854
rect 574782 60618 574866 60854
rect 575102 60618 575134 60854
rect 574514 25174 575134 60618
rect 574514 24938 574546 25174
rect 574782 24938 574866 25174
rect 575102 24938 575134 25174
rect 574514 24854 575134 24938
rect 574514 24618 574546 24854
rect 574782 24618 574866 24854
rect 575102 24618 575134 24854
rect 574514 -3226 575134 24618
rect 574514 -3462 574546 -3226
rect 574782 -3462 574866 -3226
rect 575102 -3462 575134 -3226
rect 574514 -3546 575134 -3462
rect 574514 -3782 574546 -3546
rect 574782 -3782 574866 -3546
rect 575102 -3782 575134 -3546
rect 574514 -3814 575134 -3782
rect 578234 676894 578854 709082
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 578234 676658 578266 676894
rect 578502 676658 578586 676894
rect 578822 676658 578854 676894
rect 578234 676574 578854 676658
rect 578234 676338 578266 676574
rect 578502 676338 578586 676574
rect 578822 676338 578854 676574
rect 578234 640894 578854 676338
rect 578234 640658 578266 640894
rect 578502 640658 578586 640894
rect 578822 640658 578854 640894
rect 578234 640574 578854 640658
rect 578234 640338 578266 640574
rect 578502 640338 578586 640574
rect 578822 640338 578854 640574
rect 578234 604894 578854 640338
rect 578234 604658 578266 604894
rect 578502 604658 578586 604894
rect 578822 604658 578854 604894
rect 578234 604574 578854 604658
rect 578234 604338 578266 604574
rect 578502 604338 578586 604574
rect 578822 604338 578854 604574
rect 578234 568894 578854 604338
rect 578234 568658 578266 568894
rect 578502 568658 578586 568894
rect 578822 568658 578854 568894
rect 578234 568574 578854 568658
rect 578234 568338 578266 568574
rect 578502 568338 578586 568574
rect 578822 568338 578854 568574
rect 578234 532894 578854 568338
rect 578234 532658 578266 532894
rect 578502 532658 578586 532894
rect 578822 532658 578854 532894
rect 578234 532574 578854 532658
rect 578234 532338 578266 532574
rect 578502 532338 578586 532574
rect 578822 532338 578854 532574
rect 578234 496894 578854 532338
rect 578234 496658 578266 496894
rect 578502 496658 578586 496894
rect 578822 496658 578854 496894
rect 578234 496574 578854 496658
rect 578234 496338 578266 496574
rect 578502 496338 578586 496574
rect 578822 496338 578854 496574
rect 578234 460894 578854 496338
rect 578234 460658 578266 460894
rect 578502 460658 578586 460894
rect 578822 460658 578854 460894
rect 578234 460574 578854 460658
rect 578234 460338 578266 460574
rect 578502 460338 578586 460574
rect 578822 460338 578854 460574
rect 578234 424894 578854 460338
rect 578234 424658 578266 424894
rect 578502 424658 578586 424894
rect 578822 424658 578854 424894
rect 578234 424574 578854 424658
rect 578234 424338 578266 424574
rect 578502 424338 578586 424574
rect 578822 424338 578854 424574
rect 578234 388894 578854 424338
rect 578234 388658 578266 388894
rect 578502 388658 578586 388894
rect 578822 388658 578854 388894
rect 578234 388574 578854 388658
rect 578234 388338 578266 388574
rect 578502 388338 578586 388574
rect 578822 388338 578854 388574
rect 578234 352894 578854 388338
rect 578234 352658 578266 352894
rect 578502 352658 578586 352894
rect 578822 352658 578854 352894
rect 578234 352574 578854 352658
rect 578234 352338 578266 352574
rect 578502 352338 578586 352574
rect 578822 352338 578854 352574
rect 578234 316894 578854 352338
rect 578234 316658 578266 316894
rect 578502 316658 578586 316894
rect 578822 316658 578854 316894
rect 578234 316574 578854 316658
rect 578234 316338 578266 316574
rect 578502 316338 578586 316574
rect 578822 316338 578854 316574
rect 578234 280894 578854 316338
rect 578234 280658 578266 280894
rect 578502 280658 578586 280894
rect 578822 280658 578854 280894
rect 578234 280574 578854 280658
rect 578234 280338 578266 280574
rect 578502 280338 578586 280574
rect 578822 280338 578854 280574
rect 578234 244894 578854 280338
rect 578234 244658 578266 244894
rect 578502 244658 578586 244894
rect 578822 244658 578854 244894
rect 578234 244574 578854 244658
rect 578234 244338 578266 244574
rect 578502 244338 578586 244574
rect 578822 244338 578854 244574
rect 578234 208894 578854 244338
rect 578234 208658 578266 208894
rect 578502 208658 578586 208894
rect 578822 208658 578854 208894
rect 578234 208574 578854 208658
rect 578234 208338 578266 208574
rect 578502 208338 578586 208574
rect 578822 208338 578854 208574
rect 578234 172894 578854 208338
rect 578234 172658 578266 172894
rect 578502 172658 578586 172894
rect 578822 172658 578854 172894
rect 578234 172574 578854 172658
rect 578234 172338 578266 172574
rect 578502 172338 578586 172574
rect 578822 172338 578854 172574
rect 578234 136894 578854 172338
rect 578234 136658 578266 136894
rect 578502 136658 578586 136894
rect 578822 136658 578854 136894
rect 578234 136574 578854 136658
rect 578234 136338 578266 136574
rect 578502 136338 578586 136574
rect 578822 136338 578854 136574
rect 578234 100894 578854 136338
rect 578234 100658 578266 100894
rect 578502 100658 578586 100894
rect 578822 100658 578854 100894
rect 578234 100574 578854 100658
rect 578234 100338 578266 100574
rect 578502 100338 578586 100574
rect 578822 100338 578854 100574
rect 578234 64894 578854 100338
rect 578234 64658 578266 64894
rect 578502 64658 578586 64894
rect 578822 64658 578854 64894
rect 578234 64574 578854 64658
rect 578234 64338 578266 64574
rect 578502 64338 578586 64574
rect 578822 64338 578854 64574
rect 578234 28894 578854 64338
rect 578234 28658 578266 28894
rect 578502 28658 578586 28894
rect 578822 28658 578854 28894
rect 578234 28574 578854 28658
rect 578234 28338 578266 28574
rect 578502 28338 578586 28574
rect 578822 28338 578854 28574
rect 578234 -5146 578854 28338
rect 580794 704838 581414 705830
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 580794 704602 580826 704838
rect 581062 704602 581146 704838
rect 581382 704602 581414 704838
rect 580794 704518 581414 704602
rect 580794 704282 580826 704518
rect 581062 704282 581146 704518
rect 581382 704282 581414 704518
rect 580794 687454 581414 704282
rect 580794 687218 580826 687454
rect 581062 687218 581146 687454
rect 581382 687218 581414 687454
rect 580794 687134 581414 687218
rect 580794 686898 580826 687134
rect 581062 686898 581146 687134
rect 581382 686898 581414 687134
rect 580794 651454 581414 686898
rect 580794 651218 580826 651454
rect 581062 651218 581146 651454
rect 581382 651218 581414 651454
rect 580794 651134 581414 651218
rect 580794 650898 580826 651134
rect 581062 650898 581146 651134
rect 581382 650898 581414 651134
rect 580794 615454 581414 650898
rect 580794 615218 580826 615454
rect 581062 615218 581146 615454
rect 581382 615218 581414 615454
rect 580794 615134 581414 615218
rect 580794 614898 580826 615134
rect 581062 614898 581146 615134
rect 581382 614898 581414 615134
rect 580794 579454 581414 614898
rect 580794 579218 580826 579454
rect 581062 579218 581146 579454
rect 581382 579218 581414 579454
rect 580794 579134 581414 579218
rect 580794 578898 580826 579134
rect 581062 578898 581146 579134
rect 581382 578898 581414 579134
rect 580794 543454 581414 578898
rect 580794 543218 580826 543454
rect 581062 543218 581146 543454
rect 581382 543218 581414 543454
rect 580794 543134 581414 543218
rect 580794 542898 580826 543134
rect 581062 542898 581146 543134
rect 581382 542898 581414 543134
rect 580794 507454 581414 542898
rect 580794 507218 580826 507454
rect 581062 507218 581146 507454
rect 581382 507218 581414 507454
rect 580794 507134 581414 507218
rect 580794 506898 580826 507134
rect 581062 506898 581146 507134
rect 581382 506898 581414 507134
rect 580794 471454 581414 506898
rect 580794 471218 580826 471454
rect 581062 471218 581146 471454
rect 581382 471218 581414 471454
rect 580794 471134 581414 471218
rect 580794 470898 580826 471134
rect 581062 470898 581146 471134
rect 581382 470898 581414 471134
rect 580794 435454 581414 470898
rect 580794 435218 580826 435454
rect 581062 435218 581146 435454
rect 581382 435218 581414 435454
rect 580794 435134 581414 435218
rect 580794 434898 580826 435134
rect 581062 434898 581146 435134
rect 581382 434898 581414 435134
rect 580794 399454 581414 434898
rect 580794 399218 580826 399454
rect 581062 399218 581146 399454
rect 581382 399218 581414 399454
rect 580794 399134 581414 399218
rect 580794 398898 580826 399134
rect 581062 398898 581146 399134
rect 581382 398898 581414 399134
rect 580794 363454 581414 398898
rect 580794 363218 580826 363454
rect 581062 363218 581146 363454
rect 581382 363218 581414 363454
rect 580794 363134 581414 363218
rect 580794 362898 580826 363134
rect 581062 362898 581146 363134
rect 581382 362898 581414 363134
rect 580794 327454 581414 362898
rect 580794 327218 580826 327454
rect 581062 327218 581146 327454
rect 581382 327218 581414 327454
rect 580794 327134 581414 327218
rect 580794 326898 580826 327134
rect 581062 326898 581146 327134
rect 581382 326898 581414 327134
rect 580794 291454 581414 326898
rect 580794 291218 580826 291454
rect 581062 291218 581146 291454
rect 581382 291218 581414 291454
rect 580794 291134 581414 291218
rect 580794 290898 580826 291134
rect 581062 290898 581146 291134
rect 581382 290898 581414 291134
rect 580794 255454 581414 290898
rect 580794 255218 580826 255454
rect 581062 255218 581146 255454
rect 581382 255218 581414 255454
rect 580794 255134 581414 255218
rect 580794 254898 580826 255134
rect 581062 254898 581146 255134
rect 581382 254898 581414 255134
rect 580794 219454 581414 254898
rect 580794 219218 580826 219454
rect 581062 219218 581146 219454
rect 581382 219218 581414 219454
rect 580794 219134 581414 219218
rect 580794 218898 580826 219134
rect 581062 218898 581146 219134
rect 581382 218898 581414 219134
rect 580794 183454 581414 218898
rect 580794 183218 580826 183454
rect 581062 183218 581146 183454
rect 581382 183218 581414 183454
rect 580794 183134 581414 183218
rect 580794 182898 580826 183134
rect 581062 182898 581146 183134
rect 581382 182898 581414 183134
rect 580794 147454 581414 182898
rect 580794 147218 580826 147454
rect 581062 147218 581146 147454
rect 581382 147218 581414 147454
rect 580794 147134 581414 147218
rect 580794 146898 580826 147134
rect 581062 146898 581146 147134
rect 581382 146898 581414 147134
rect 580794 111454 581414 146898
rect 580794 111218 580826 111454
rect 581062 111218 581146 111454
rect 581382 111218 581414 111454
rect 580794 111134 581414 111218
rect 580794 110898 580826 111134
rect 581062 110898 581146 111134
rect 581382 110898 581414 111134
rect 580794 75454 581414 110898
rect 580794 75218 580826 75454
rect 581062 75218 581146 75454
rect 581382 75218 581414 75454
rect 580794 75134 581414 75218
rect 580794 74898 580826 75134
rect 581062 74898 581146 75134
rect 581382 74898 581414 75134
rect 580794 39454 581414 74898
rect 580794 39218 580826 39454
rect 581062 39218 581146 39454
rect 581382 39218 581414 39454
rect 580794 39134 581414 39218
rect 580794 38898 580826 39134
rect 581062 38898 581146 39134
rect 581382 38898 581414 39134
rect 580794 3454 581414 38898
rect 580794 3218 580826 3454
rect 581062 3218 581146 3454
rect 581382 3218 581414 3454
rect 580794 3134 581414 3218
rect 580794 2898 580826 3134
rect 581062 2898 581146 3134
rect 581382 2898 581414 3134
rect 580794 -346 581414 2898
rect 580794 -582 580826 -346
rect 581062 -582 581146 -346
rect 581382 -582 581414 -346
rect 580794 -666 581414 -582
rect 580794 -902 580826 -666
rect 581062 -902 581146 -666
rect 581382 -902 581414 -666
rect 580794 -1894 581414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 578234 -5382 578266 -5146
rect 578502 -5382 578586 -5146
rect 578822 -5382 578854 -5146
rect 578234 -5466 578854 -5382
rect 578234 -5702 578266 -5466
rect 578502 -5702 578586 -5466
rect 578822 -5702 578854 -5466
rect 578234 -5734 578854 -5702
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 571954 -6342 571986 -6106
rect 572222 -6342 572306 -6106
rect 572542 -6342 572574 -6106
rect 571954 -6426 572574 -6342
rect 571954 -6662 571986 -6426
rect 572222 -6662 572306 -6426
rect 572542 -6662 572574 -6426
rect 571954 -7654 572574 -6662
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 11986 710362 12222 710598
rect 12306 710362 12542 710598
rect 11986 710042 12222 710278
rect 12306 710042 12542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 8266 708442 8502 708678
rect 8586 708442 8822 708678
rect 8266 708122 8502 708358
rect 8586 708122 8822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 4546 706522 4782 706758
rect 4866 706522 5102 706758
rect 4546 706202 4782 706438
rect 4866 706202 5102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 826 704602 1062 704838
rect 1146 704602 1382 704838
rect 826 704282 1062 704518
rect 1146 704282 1382 704518
rect 826 687218 1062 687454
rect 1146 687218 1382 687454
rect 826 686898 1062 687134
rect 1146 686898 1382 687134
rect 826 651218 1062 651454
rect 1146 651218 1382 651454
rect 826 650898 1062 651134
rect 1146 650898 1382 651134
rect 826 615218 1062 615454
rect 1146 615218 1382 615454
rect 826 614898 1062 615134
rect 1146 614898 1382 615134
rect 826 579218 1062 579454
rect 1146 579218 1382 579454
rect 826 578898 1062 579134
rect 1146 578898 1382 579134
rect 826 543218 1062 543454
rect 1146 543218 1382 543454
rect 826 542898 1062 543134
rect 1146 542898 1382 543134
rect 826 507218 1062 507454
rect 1146 507218 1382 507454
rect 826 506898 1062 507134
rect 1146 506898 1382 507134
rect 826 471218 1062 471454
rect 1146 471218 1382 471454
rect 826 470898 1062 471134
rect 1146 470898 1382 471134
rect 826 435218 1062 435454
rect 1146 435218 1382 435454
rect 826 434898 1062 435134
rect 1146 434898 1382 435134
rect 826 399218 1062 399454
rect 1146 399218 1382 399454
rect 826 398898 1062 399134
rect 1146 398898 1382 399134
rect 826 363218 1062 363454
rect 1146 363218 1382 363454
rect 826 362898 1062 363134
rect 1146 362898 1382 363134
rect 826 327218 1062 327454
rect 1146 327218 1382 327454
rect 826 326898 1062 327134
rect 1146 326898 1382 327134
rect 826 291218 1062 291454
rect 1146 291218 1382 291454
rect 826 290898 1062 291134
rect 1146 290898 1382 291134
rect 826 255218 1062 255454
rect 1146 255218 1382 255454
rect 826 254898 1062 255134
rect 1146 254898 1382 255134
rect 826 219218 1062 219454
rect 1146 219218 1382 219454
rect 826 218898 1062 219134
rect 1146 218898 1382 219134
rect 826 183218 1062 183454
rect 1146 183218 1382 183454
rect 826 182898 1062 183134
rect 1146 182898 1382 183134
rect 826 147218 1062 147454
rect 1146 147218 1382 147454
rect 826 146898 1062 147134
rect 1146 146898 1382 147134
rect 826 111218 1062 111454
rect 1146 111218 1382 111454
rect 826 110898 1062 111134
rect 1146 110898 1382 111134
rect 826 75218 1062 75454
rect 1146 75218 1382 75454
rect 826 74898 1062 75134
rect 1146 74898 1382 75134
rect 826 39218 1062 39454
rect 1146 39218 1382 39454
rect 826 38898 1062 39134
rect 1146 38898 1382 39134
rect 826 3218 1062 3454
rect 1146 3218 1382 3454
rect 826 2898 1062 3134
rect 1146 2898 1382 3134
rect 826 -582 1062 -346
rect 1146 -582 1382 -346
rect 826 -902 1062 -666
rect 1146 -902 1382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 4546 690938 4782 691174
rect 4866 690938 5102 691174
rect 4546 690618 4782 690854
rect 4866 690618 5102 690854
rect 4546 654938 4782 655174
rect 4866 654938 5102 655174
rect 4546 654618 4782 654854
rect 4866 654618 5102 654854
rect 4546 618938 4782 619174
rect 4866 618938 5102 619174
rect 4546 618618 4782 618854
rect 4866 618618 5102 618854
rect 4546 582938 4782 583174
rect 4866 582938 5102 583174
rect 4546 582618 4782 582854
rect 4866 582618 5102 582854
rect 4546 546938 4782 547174
rect 4866 546938 5102 547174
rect 4546 546618 4782 546854
rect 4866 546618 5102 546854
rect 4546 510938 4782 511174
rect 4866 510938 5102 511174
rect 4546 510618 4782 510854
rect 4866 510618 5102 510854
rect 4546 474938 4782 475174
rect 4866 474938 5102 475174
rect 4546 474618 4782 474854
rect 4866 474618 5102 474854
rect 4546 438938 4782 439174
rect 4866 438938 5102 439174
rect 4546 438618 4782 438854
rect 4866 438618 5102 438854
rect 4546 402938 4782 403174
rect 4866 402938 5102 403174
rect 4546 402618 4782 402854
rect 4866 402618 5102 402854
rect 4546 366938 4782 367174
rect 4866 366938 5102 367174
rect 4546 366618 4782 366854
rect 4866 366618 5102 366854
rect 4546 330938 4782 331174
rect 4866 330938 5102 331174
rect 4546 330618 4782 330854
rect 4866 330618 5102 330854
rect 4546 294938 4782 295174
rect 4866 294938 5102 295174
rect 4546 294618 4782 294854
rect 4866 294618 5102 294854
rect 4546 258938 4782 259174
rect 4866 258938 5102 259174
rect 4546 258618 4782 258854
rect 4866 258618 5102 258854
rect 4546 222938 4782 223174
rect 4866 222938 5102 223174
rect 4546 222618 4782 222854
rect 4866 222618 5102 222854
rect 4546 186938 4782 187174
rect 4866 186938 5102 187174
rect 4546 186618 4782 186854
rect 4866 186618 5102 186854
rect 4546 150938 4782 151174
rect 4866 150938 5102 151174
rect 4546 150618 4782 150854
rect 4866 150618 5102 150854
rect 4546 114938 4782 115174
rect 4866 114938 5102 115174
rect 4546 114618 4782 114854
rect 4866 114618 5102 114854
rect 4546 78938 4782 79174
rect 4866 78938 5102 79174
rect 4546 78618 4782 78854
rect 4866 78618 5102 78854
rect 4546 42938 4782 43174
rect 4866 42938 5102 43174
rect 4546 42618 4782 42854
rect 4866 42618 5102 42854
rect 4546 6938 4782 7174
rect 4866 6938 5102 7174
rect 4546 6618 4782 6854
rect 4866 6618 5102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 4546 -2502 4782 -2266
rect 4866 -2502 5102 -2266
rect 4546 -2822 4782 -2586
rect 4866 -2822 5102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 8266 694658 8502 694894
rect 8586 694658 8822 694894
rect 8266 694338 8502 694574
rect 8586 694338 8822 694574
rect 8266 658658 8502 658894
rect 8586 658658 8822 658894
rect 8266 658338 8502 658574
rect 8586 658338 8822 658574
rect 8266 622658 8502 622894
rect 8586 622658 8822 622894
rect 8266 622338 8502 622574
rect 8586 622338 8822 622574
rect 8266 586658 8502 586894
rect 8586 586658 8822 586894
rect 8266 586338 8502 586574
rect 8586 586338 8822 586574
rect 8266 550658 8502 550894
rect 8586 550658 8822 550894
rect 8266 550338 8502 550574
rect 8586 550338 8822 550574
rect 8266 514658 8502 514894
rect 8586 514658 8822 514894
rect 8266 514338 8502 514574
rect 8586 514338 8822 514574
rect 8266 478658 8502 478894
rect 8586 478658 8822 478894
rect 8266 478338 8502 478574
rect 8586 478338 8822 478574
rect 8266 442658 8502 442894
rect 8586 442658 8822 442894
rect 8266 442338 8502 442574
rect 8586 442338 8822 442574
rect 8266 406658 8502 406894
rect 8586 406658 8822 406894
rect 8266 406338 8502 406574
rect 8586 406338 8822 406574
rect 8266 370658 8502 370894
rect 8586 370658 8822 370894
rect 8266 370338 8502 370574
rect 8586 370338 8822 370574
rect 8266 334658 8502 334894
rect 8586 334658 8822 334894
rect 8266 334338 8502 334574
rect 8586 334338 8822 334574
rect 8266 298658 8502 298894
rect 8586 298658 8822 298894
rect 8266 298338 8502 298574
rect 8586 298338 8822 298574
rect 8266 262658 8502 262894
rect 8586 262658 8822 262894
rect 8266 262338 8502 262574
rect 8586 262338 8822 262574
rect 8266 226658 8502 226894
rect 8586 226658 8822 226894
rect 8266 226338 8502 226574
rect 8586 226338 8822 226574
rect 8266 190658 8502 190894
rect 8586 190658 8822 190894
rect 8266 190338 8502 190574
rect 8586 190338 8822 190574
rect 8266 154658 8502 154894
rect 8586 154658 8822 154894
rect 8266 154338 8502 154574
rect 8586 154338 8822 154574
rect 8266 118658 8502 118894
rect 8586 118658 8822 118894
rect 8266 118338 8502 118574
rect 8586 118338 8822 118574
rect 8266 82658 8502 82894
rect 8586 82658 8822 82894
rect 8266 82338 8502 82574
rect 8586 82338 8822 82574
rect 8266 46658 8502 46894
rect 8586 46658 8822 46894
rect 8266 46338 8502 46574
rect 8586 46338 8822 46574
rect 8266 10658 8502 10894
rect 8586 10658 8822 10894
rect 8266 10338 8502 10574
rect 8586 10338 8822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 10826 705562 11062 705798
rect 11146 705562 11382 705798
rect 10826 705242 11062 705478
rect 11146 705242 11382 705478
rect 10826 669218 11062 669454
rect 11146 669218 11382 669454
rect 10826 668898 11062 669134
rect 11146 668898 11382 669134
rect 10826 633218 11062 633454
rect 11146 633218 11382 633454
rect 10826 632898 11062 633134
rect 11146 632898 11382 633134
rect 10826 597218 11062 597454
rect 11146 597218 11382 597454
rect 10826 596898 11062 597134
rect 11146 596898 11382 597134
rect 10826 561218 11062 561454
rect 11146 561218 11382 561454
rect 10826 560898 11062 561134
rect 11146 560898 11382 561134
rect 10826 525218 11062 525454
rect 11146 525218 11382 525454
rect 10826 524898 11062 525134
rect 11146 524898 11382 525134
rect 10826 489218 11062 489454
rect 11146 489218 11382 489454
rect 10826 488898 11062 489134
rect 11146 488898 11382 489134
rect 10826 453218 11062 453454
rect 11146 453218 11382 453454
rect 10826 452898 11062 453134
rect 11146 452898 11382 453134
rect 10826 417218 11062 417454
rect 11146 417218 11382 417454
rect 10826 416898 11062 417134
rect 11146 416898 11382 417134
rect 10826 381218 11062 381454
rect 11146 381218 11382 381454
rect 10826 380898 11062 381134
rect 11146 380898 11382 381134
rect 10826 345218 11062 345454
rect 11146 345218 11382 345454
rect 10826 344898 11062 345134
rect 11146 344898 11382 345134
rect 10826 309218 11062 309454
rect 11146 309218 11382 309454
rect 10826 308898 11062 309134
rect 11146 308898 11382 309134
rect 10826 273218 11062 273454
rect 11146 273218 11382 273454
rect 10826 272898 11062 273134
rect 11146 272898 11382 273134
rect 10826 237218 11062 237454
rect 11146 237218 11382 237454
rect 10826 236898 11062 237134
rect 11146 236898 11382 237134
rect 10826 201218 11062 201454
rect 11146 201218 11382 201454
rect 10826 200898 11062 201134
rect 11146 200898 11382 201134
rect 10826 165218 11062 165454
rect 11146 165218 11382 165454
rect 10826 164898 11062 165134
rect 11146 164898 11382 165134
rect 10826 129218 11062 129454
rect 11146 129218 11382 129454
rect 10826 128898 11062 129134
rect 11146 128898 11382 129134
rect 10826 93218 11062 93454
rect 11146 93218 11382 93454
rect 10826 92898 11062 93134
rect 11146 92898 11382 93134
rect 10826 57218 11062 57454
rect 11146 57218 11382 57454
rect 10826 56898 11062 57134
rect 11146 56898 11382 57134
rect 10826 21218 11062 21454
rect 11146 21218 11382 21454
rect 10826 20898 11062 21134
rect 11146 20898 11382 21134
rect 10826 -1542 11062 -1306
rect 11146 -1542 11382 -1306
rect 10826 -1862 11062 -1626
rect 11146 -1862 11382 -1626
rect 21986 711322 22222 711558
rect 22306 711322 22542 711558
rect 21986 711002 22222 711238
rect 22306 711002 22542 711238
rect 18266 709402 18502 709638
rect 18586 709402 18822 709638
rect 18266 709082 18502 709318
rect 18586 709082 18822 709318
rect 11986 698378 12222 698614
rect 12306 698378 12542 698614
rect 11986 698058 12222 698294
rect 12306 698058 12542 698294
rect 11986 662378 12222 662614
rect 12306 662378 12542 662614
rect 11986 662058 12222 662294
rect 12306 662058 12542 662294
rect 11986 626378 12222 626614
rect 12306 626378 12542 626614
rect 11986 626058 12222 626294
rect 12306 626058 12542 626294
rect 11986 590378 12222 590614
rect 12306 590378 12542 590614
rect 11986 590058 12222 590294
rect 12306 590058 12542 590294
rect 11986 554378 12222 554614
rect 12306 554378 12542 554614
rect 11986 554058 12222 554294
rect 12306 554058 12542 554294
rect 11986 518378 12222 518614
rect 12306 518378 12542 518614
rect 11986 518058 12222 518294
rect 12306 518058 12542 518294
rect 11986 482378 12222 482614
rect 12306 482378 12542 482614
rect 11986 482058 12222 482294
rect 12306 482058 12542 482294
rect 11986 446378 12222 446614
rect 12306 446378 12542 446614
rect 11986 446058 12222 446294
rect 12306 446058 12542 446294
rect 11986 410378 12222 410614
rect 12306 410378 12542 410614
rect 11986 410058 12222 410294
rect 12306 410058 12542 410294
rect 11986 374378 12222 374614
rect 12306 374378 12542 374614
rect 11986 374058 12222 374294
rect 12306 374058 12542 374294
rect 11986 338378 12222 338614
rect 12306 338378 12542 338614
rect 11986 338058 12222 338294
rect 12306 338058 12542 338294
rect 11986 302378 12222 302614
rect 12306 302378 12542 302614
rect 11986 302058 12222 302294
rect 12306 302058 12542 302294
rect 11986 266378 12222 266614
rect 12306 266378 12542 266614
rect 11986 266058 12222 266294
rect 12306 266058 12542 266294
rect 11986 230378 12222 230614
rect 12306 230378 12542 230614
rect 11986 230058 12222 230294
rect 12306 230058 12542 230294
rect 11986 194378 12222 194614
rect 12306 194378 12542 194614
rect 11986 194058 12222 194294
rect 12306 194058 12542 194294
rect 11986 158378 12222 158614
rect 12306 158378 12542 158614
rect 11986 158058 12222 158294
rect 12306 158058 12542 158294
rect 11986 122378 12222 122614
rect 12306 122378 12542 122614
rect 11986 122058 12222 122294
rect 12306 122058 12542 122294
rect 11986 86378 12222 86614
rect 12306 86378 12542 86614
rect 11986 86058 12222 86294
rect 12306 86058 12542 86294
rect 11986 50378 12222 50614
rect 12306 50378 12542 50614
rect 11986 50058 12222 50294
rect 12306 50058 12542 50294
rect 11986 14378 12222 14614
rect 12306 14378 12542 14614
rect 11986 14058 12222 14294
rect 12306 14058 12542 14294
rect 8266 -4422 8502 -4186
rect 8586 -4422 8822 -4186
rect 8266 -4742 8502 -4506
rect 8586 -4742 8822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 14546 707482 14782 707718
rect 14866 707482 15102 707718
rect 14546 707162 14782 707398
rect 14866 707162 15102 707398
rect 14546 672938 14782 673174
rect 14866 672938 15102 673174
rect 14546 672618 14782 672854
rect 14866 672618 15102 672854
rect 14546 636938 14782 637174
rect 14866 636938 15102 637174
rect 14546 636618 14782 636854
rect 14866 636618 15102 636854
rect 14546 600938 14782 601174
rect 14866 600938 15102 601174
rect 14546 600618 14782 600854
rect 14866 600618 15102 600854
rect 14546 564938 14782 565174
rect 14866 564938 15102 565174
rect 14546 564618 14782 564854
rect 14866 564618 15102 564854
rect 14546 528938 14782 529174
rect 14866 528938 15102 529174
rect 14546 528618 14782 528854
rect 14866 528618 15102 528854
rect 14546 492938 14782 493174
rect 14866 492938 15102 493174
rect 14546 492618 14782 492854
rect 14866 492618 15102 492854
rect 14546 456938 14782 457174
rect 14866 456938 15102 457174
rect 14546 456618 14782 456854
rect 14866 456618 15102 456854
rect 14546 420938 14782 421174
rect 14866 420938 15102 421174
rect 14546 420618 14782 420854
rect 14866 420618 15102 420854
rect 14546 384938 14782 385174
rect 14866 384938 15102 385174
rect 14546 384618 14782 384854
rect 14866 384618 15102 384854
rect 14546 348938 14782 349174
rect 14866 348938 15102 349174
rect 14546 348618 14782 348854
rect 14866 348618 15102 348854
rect 14546 312938 14782 313174
rect 14866 312938 15102 313174
rect 14546 312618 14782 312854
rect 14866 312618 15102 312854
rect 14546 276938 14782 277174
rect 14866 276938 15102 277174
rect 14546 276618 14782 276854
rect 14866 276618 15102 276854
rect 14546 240938 14782 241174
rect 14866 240938 15102 241174
rect 14546 240618 14782 240854
rect 14866 240618 15102 240854
rect 14546 204938 14782 205174
rect 14866 204938 15102 205174
rect 14546 204618 14782 204854
rect 14866 204618 15102 204854
rect 14546 168938 14782 169174
rect 14866 168938 15102 169174
rect 14546 168618 14782 168854
rect 14866 168618 15102 168854
rect 14546 132938 14782 133174
rect 14866 132938 15102 133174
rect 14546 132618 14782 132854
rect 14866 132618 15102 132854
rect 14546 96938 14782 97174
rect 14866 96938 15102 97174
rect 14546 96618 14782 96854
rect 14866 96618 15102 96854
rect 18266 676658 18502 676894
rect 18586 676658 18822 676894
rect 18266 676338 18502 676574
rect 18586 676338 18822 676574
rect 18266 640658 18502 640894
rect 18586 640658 18822 640894
rect 18266 640338 18502 640574
rect 18586 640338 18822 640574
rect 18266 604658 18502 604894
rect 18586 604658 18822 604894
rect 18266 604338 18502 604574
rect 18586 604338 18822 604574
rect 18266 568658 18502 568894
rect 18586 568658 18822 568894
rect 18266 568338 18502 568574
rect 18586 568338 18822 568574
rect 18266 532658 18502 532894
rect 18586 532658 18822 532894
rect 18266 532338 18502 532574
rect 18586 532338 18822 532574
rect 18266 496658 18502 496894
rect 18586 496658 18822 496894
rect 18266 496338 18502 496574
rect 18586 496338 18822 496574
rect 18266 460658 18502 460894
rect 18586 460658 18822 460894
rect 18266 460338 18502 460574
rect 18586 460338 18822 460574
rect 18266 424658 18502 424894
rect 18586 424658 18822 424894
rect 18266 424338 18502 424574
rect 18586 424338 18822 424574
rect 18266 388658 18502 388894
rect 18586 388658 18822 388894
rect 18266 388338 18502 388574
rect 18586 388338 18822 388574
rect 18266 352658 18502 352894
rect 18586 352658 18822 352894
rect 18266 352338 18502 352574
rect 18586 352338 18822 352574
rect 18266 316658 18502 316894
rect 18586 316658 18822 316894
rect 18266 316338 18502 316574
rect 18586 316338 18822 316574
rect 18266 280658 18502 280894
rect 18586 280658 18822 280894
rect 18266 280338 18502 280574
rect 18586 280338 18822 280574
rect 18266 244658 18502 244894
rect 18586 244658 18822 244894
rect 18266 244338 18502 244574
rect 18586 244338 18822 244574
rect 18266 208658 18502 208894
rect 18586 208658 18822 208894
rect 18266 208338 18502 208574
rect 18586 208338 18822 208574
rect 18266 172658 18502 172894
rect 18586 172658 18822 172894
rect 18266 172338 18502 172574
rect 18586 172338 18822 172574
rect 18266 136658 18502 136894
rect 18586 136658 18822 136894
rect 18266 136338 18502 136574
rect 18586 136338 18822 136574
rect 18266 100658 18502 100894
rect 18586 100658 18822 100894
rect 18266 100338 18502 100574
rect 18586 100338 18822 100574
rect 20826 704602 21062 704838
rect 21146 704602 21382 704838
rect 20826 704282 21062 704518
rect 21146 704282 21382 704518
rect 20826 687218 21062 687454
rect 21146 687218 21382 687454
rect 20826 686898 21062 687134
rect 21146 686898 21382 687134
rect 20826 651218 21062 651454
rect 21146 651218 21382 651454
rect 20826 650898 21062 651134
rect 21146 650898 21382 651134
rect 20826 615218 21062 615454
rect 21146 615218 21382 615454
rect 20826 614898 21062 615134
rect 21146 614898 21382 615134
rect 20826 579218 21062 579454
rect 21146 579218 21382 579454
rect 20826 578898 21062 579134
rect 21146 578898 21382 579134
rect 20826 543218 21062 543454
rect 21146 543218 21382 543454
rect 20826 542898 21062 543134
rect 21146 542898 21382 543134
rect 20826 507218 21062 507454
rect 21146 507218 21382 507454
rect 20826 506898 21062 507134
rect 21146 506898 21382 507134
rect 20826 471218 21062 471454
rect 21146 471218 21382 471454
rect 20826 470898 21062 471134
rect 21146 470898 21382 471134
rect 20826 435218 21062 435454
rect 21146 435218 21382 435454
rect 20826 434898 21062 435134
rect 21146 434898 21382 435134
rect 20826 399218 21062 399454
rect 21146 399218 21382 399454
rect 20826 398898 21062 399134
rect 21146 398898 21382 399134
rect 20826 363218 21062 363454
rect 21146 363218 21382 363454
rect 20826 362898 21062 363134
rect 21146 362898 21382 363134
rect 20826 327218 21062 327454
rect 21146 327218 21382 327454
rect 20826 326898 21062 327134
rect 21146 326898 21382 327134
rect 20826 291218 21062 291454
rect 21146 291218 21382 291454
rect 20826 290898 21062 291134
rect 21146 290898 21382 291134
rect 20826 255218 21062 255454
rect 21146 255218 21382 255454
rect 20826 254898 21062 255134
rect 21146 254898 21382 255134
rect 20826 219218 21062 219454
rect 21146 219218 21382 219454
rect 20826 218898 21062 219134
rect 21146 218898 21382 219134
rect 20826 183218 21062 183454
rect 21146 183218 21382 183454
rect 20826 182898 21062 183134
rect 21146 182898 21382 183134
rect 20826 147218 21062 147454
rect 21146 147218 21382 147454
rect 20826 146898 21062 147134
rect 21146 146898 21382 147134
rect 20826 111218 21062 111454
rect 21146 111218 21382 111454
rect 20826 110898 21062 111134
rect 21146 110898 21382 111134
rect 20826 75218 21062 75454
rect 21146 75218 21382 75454
rect 20826 74898 21062 75134
rect 21146 74898 21382 75134
rect 31986 710362 32222 710598
rect 32306 710362 32542 710598
rect 31986 710042 32222 710278
rect 32306 710042 32542 710278
rect 28266 708442 28502 708678
rect 28586 708442 28822 708678
rect 28266 708122 28502 708358
rect 28586 708122 28822 708358
rect 21986 680378 22222 680614
rect 22306 680378 22542 680614
rect 21986 680058 22222 680294
rect 22306 680058 22542 680294
rect 21986 644378 22222 644614
rect 22306 644378 22542 644614
rect 21986 644058 22222 644294
rect 22306 644058 22542 644294
rect 21986 608378 22222 608614
rect 22306 608378 22542 608614
rect 21986 608058 22222 608294
rect 22306 608058 22542 608294
rect 21986 572378 22222 572614
rect 22306 572378 22542 572614
rect 21986 572058 22222 572294
rect 22306 572058 22542 572294
rect 21986 536378 22222 536614
rect 22306 536378 22542 536614
rect 21986 536058 22222 536294
rect 22306 536058 22542 536294
rect 21986 500378 22222 500614
rect 22306 500378 22542 500614
rect 21986 500058 22222 500294
rect 22306 500058 22542 500294
rect 21986 464378 22222 464614
rect 22306 464378 22542 464614
rect 21986 464058 22222 464294
rect 22306 464058 22542 464294
rect 21986 428378 22222 428614
rect 22306 428378 22542 428614
rect 21986 428058 22222 428294
rect 22306 428058 22542 428294
rect 21986 392378 22222 392614
rect 22306 392378 22542 392614
rect 21986 392058 22222 392294
rect 22306 392058 22542 392294
rect 21986 356378 22222 356614
rect 22306 356378 22542 356614
rect 21986 356058 22222 356294
rect 22306 356058 22542 356294
rect 21986 320378 22222 320614
rect 22306 320378 22542 320614
rect 21986 320058 22222 320294
rect 22306 320058 22542 320294
rect 21986 284378 22222 284614
rect 22306 284378 22542 284614
rect 21986 284058 22222 284294
rect 22306 284058 22542 284294
rect 21986 248378 22222 248614
rect 22306 248378 22542 248614
rect 21986 248058 22222 248294
rect 22306 248058 22542 248294
rect 21986 212378 22222 212614
rect 22306 212378 22542 212614
rect 21986 212058 22222 212294
rect 22306 212058 22542 212294
rect 21986 176378 22222 176614
rect 22306 176378 22542 176614
rect 21986 176058 22222 176294
rect 22306 176058 22542 176294
rect 21986 140378 22222 140614
rect 22306 140378 22542 140614
rect 21986 140058 22222 140294
rect 22306 140058 22542 140294
rect 21986 104378 22222 104614
rect 22306 104378 22542 104614
rect 21986 104058 22222 104294
rect 22306 104058 22542 104294
rect 24546 706522 24782 706758
rect 24866 706522 25102 706758
rect 24546 706202 24782 706438
rect 24866 706202 25102 706438
rect 24546 690938 24782 691174
rect 24866 690938 25102 691174
rect 24546 690618 24782 690854
rect 24866 690618 25102 690854
rect 24546 654938 24782 655174
rect 24866 654938 25102 655174
rect 24546 654618 24782 654854
rect 24866 654618 25102 654854
rect 24546 618938 24782 619174
rect 24866 618938 25102 619174
rect 24546 618618 24782 618854
rect 24866 618618 25102 618854
rect 24546 582938 24782 583174
rect 24866 582938 25102 583174
rect 24546 582618 24782 582854
rect 24866 582618 25102 582854
rect 24546 546938 24782 547174
rect 24866 546938 25102 547174
rect 24546 546618 24782 546854
rect 24866 546618 25102 546854
rect 24546 510938 24782 511174
rect 24866 510938 25102 511174
rect 24546 510618 24782 510854
rect 24866 510618 25102 510854
rect 24546 474938 24782 475174
rect 24866 474938 25102 475174
rect 24546 474618 24782 474854
rect 24866 474618 25102 474854
rect 24546 438938 24782 439174
rect 24866 438938 25102 439174
rect 24546 438618 24782 438854
rect 24866 438618 25102 438854
rect 24546 402938 24782 403174
rect 24866 402938 25102 403174
rect 24546 402618 24782 402854
rect 24866 402618 25102 402854
rect 24546 366938 24782 367174
rect 24866 366938 25102 367174
rect 24546 366618 24782 366854
rect 24866 366618 25102 366854
rect 24546 330938 24782 331174
rect 24866 330938 25102 331174
rect 24546 330618 24782 330854
rect 24866 330618 25102 330854
rect 24546 294938 24782 295174
rect 24866 294938 25102 295174
rect 24546 294618 24782 294854
rect 24866 294618 25102 294854
rect 24546 258938 24782 259174
rect 24866 258938 25102 259174
rect 24546 258618 24782 258854
rect 24866 258618 25102 258854
rect 24546 222938 24782 223174
rect 24866 222938 25102 223174
rect 24546 222618 24782 222854
rect 24866 222618 25102 222854
rect 24546 186938 24782 187174
rect 24866 186938 25102 187174
rect 24546 186618 24782 186854
rect 24866 186618 25102 186854
rect 24546 150938 24782 151174
rect 24866 150938 25102 151174
rect 24546 150618 24782 150854
rect 24866 150618 25102 150854
rect 24546 114938 24782 115174
rect 24866 114938 25102 115174
rect 24546 114618 24782 114854
rect 24866 114618 25102 114854
rect 24546 78938 24782 79174
rect 24866 78938 25102 79174
rect 24546 78618 24782 78854
rect 24866 78618 25102 78854
rect 28266 694658 28502 694894
rect 28586 694658 28822 694894
rect 28266 694338 28502 694574
rect 28586 694338 28822 694574
rect 28266 658658 28502 658894
rect 28586 658658 28822 658894
rect 28266 658338 28502 658574
rect 28586 658338 28822 658574
rect 28266 622658 28502 622894
rect 28586 622658 28822 622894
rect 28266 622338 28502 622574
rect 28586 622338 28822 622574
rect 28266 586658 28502 586894
rect 28586 586658 28822 586894
rect 28266 586338 28502 586574
rect 28586 586338 28822 586574
rect 28266 550658 28502 550894
rect 28586 550658 28822 550894
rect 28266 550338 28502 550574
rect 28586 550338 28822 550574
rect 28266 514658 28502 514894
rect 28586 514658 28822 514894
rect 28266 514338 28502 514574
rect 28586 514338 28822 514574
rect 28266 478658 28502 478894
rect 28586 478658 28822 478894
rect 28266 478338 28502 478574
rect 28586 478338 28822 478574
rect 28266 442658 28502 442894
rect 28586 442658 28822 442894
rect 28266 442338 28502 442574
rect 28586 442338 28822 442574
rect 28266 406658 28502 406894
rect 28586 406658 28822 406894
rect 28266 406338 28502 406574
rect 28586 406338 28822 406574
rect 28266 370658 28502 370894
rect 28586 370658 28822 370894
rect 28266 370338 28502 370574
rect 28586 370338 28822 370574
rect 28266 334658 28502 334894
rect 28586 334658 28822 334894
rect 28266 334338 28502 334574
rect 28586 334338 28822 334574
rect 28266 298658 28502 298894
rect 28586 298658 28822 298894
rect 28266 298338 28502 298574
rect 28586 298338 28822 298574
rect 28266 262658 28502 262894
rect 28586 262658 28822 262894
rect 28266 262338 28502 262574
rect 28586 262338 28822 262574
rect 28266 226658 28502 226894
rect 28586 226658 28822 226894
rect 28266 226338 28502 226574
rect 28586 226338 28822 226574
rect 28266 190658 28502 190894
rect 28586 190658 28822 190894
rect 28266 190338 28502 190574
rect 28586 190338 28822 190574
rect 28266 154658 28502 154894
rect 28586 154658 28822 154894
rect 28266 154338 28502 154574
rect 28586 154338 28822 154574
rect 28266 118658 28502 118894
rect 28586 118658 28822 118894
rect 28266 118338 28502 118574
rect 28586 118338 28822 118574
rect 28266 82658 28502 82894
rect 28586 82658 28822 82894
rect 28266 82338 28502 82574
rect 28586 82338 28822 82574
rect 30826 705562 31062 705798
rect 31146 705562 31382 705798
rect 30826 705242 31062 705478
rect 31146 705242 31382 705478
rect 30826 669218 31062 669454
rect 31146 669218 31382 669454
rect 30826 668898 31062 669134
rect 31146 668898 31382 669134
rect 30826 633218 31062 633454
rect 31146 633218 31382 633454
rect 30826 632898 31062 633134
rect 31146 632898 31382 633134
rect 30826 597218 31062 597454
rect 31146 597218 31382 597454
rect 30826 596898 31062 597134
rect 31146 596898 31382 597134
rect 30826 561218 31062 561454
rect 31146 561218 31382 561454
rect 30826 560898 31062 561134
rect 31146 560898 31382 561134
rect 30826 525218 31062 525454
rect 31146 525218 31382 525454
rect 30826 524898 31062 525134
rect 31146 524898 31382 525134
rect 30826 489218 31062 489454
rect 31146 489218 31382 489454
rect 30826 488898 31062 489134
rect 31146 488898 31382 489134
rect 30826 453218 31062 453454
rect 31146 453218 31382 453454
rect 30826 452898 31062 453134
rect 31146 452898 31382 453134
rect 30826 417218 31062 417454
rect 31146 417218 31382 417454
rect 30826 416898 31062 417134
rect 31146 416898 31382 417134
rect 30826 381218 31062 381454
rect 31146 381218 31382 381454
rect 30826 380898 31062 381134
rect 31146 380898 31382 381134
rect 30826 345218 31062 345454
rect 31146 345218 31382 345454
rect 30826 344898 31062 345134
rect 31146 344898 31382 345134
rect 30826 309218 31062 309454
rect 31146 309218 31382 309454
rect 30826 308898 31062 309134
rect 31146 308898 31382 309134
rect 30826 273218 31062 273454
rect 31146 273218 31382 273454
rect 30826 272898 31062 273134
rect 31146 272898 31382 273134
rect 30826 237218 31062 237454
rect 31146 237218 31382 237454
rect 30826 236898 31062 237134
rect 31146 236898 31382 237134
rect 30826 201218 31062 201454
rect 31146 201218 31382 201454
rect 30826 200898 31062 201134
rect 31146 200898 31382 201134
rect 30826 165218 31062 165454
rect 31146 165218 31382 165454
rect 30826 164898 31062 165134
rect 31146 164898 31382 165134
rect 30826 129218 31062 129454
rect 31146 129218 31382 129454
rect 30826 128898 31062 129134
rect 31146 128898 31382 129134
rect 30826 93218 31062 93454
rect 31146 93218 31382 93454
rect 30826 92898 31062 93134
rect 31146 92898 31382 93134
rect 41986 711322 42222 711558
rect 42306 711322 42542 711558
rect 41986 711002 42222 711238
rect 42306 711002 42542 711238
rect 38266 709402 38502 709638
rect 38586 709402 38822 709638
rect 38266 709082 38502 709318
rect 38586 709082 38822 709318
rect 31986 698378 32222 698614
rect 32306 698378 32542 698614
rect 31986 698058 32222 698294
rect 32306 698058 32542 698294
rect 31986 662378 32222 662614
rect 32306 662378 32542 662614
rect 31986 662058 32222 662294
rect 32306 662058 32542 662294
rect 31986 626378 32222 626614
rect 32306 626378 32542 626614
rect 31986 626058 32222 626294
rect 32306 626058 32542 626294
rect 31986 590378 32222 590614
rect 32306 590378 32542 590614
rect 31986 590058 32222 590294
rect 32306 590058 32542 590294
rect 31986 554378 32222 554614
rect 32306 554378 32542 554614
rect 31986 554058 32222 554294
rect 32306 554058 32542 554294
rect 31986 518378 32222 518614
rect 32306 518378 32542 518614
rect 31986 518058 32222 518294
rect 32306 518058 32542 518294
rect 31986 482378 32222 482614
rect 32306 482378 32542 482614
rect 31986 482058 32222 482294
rect 32306 482058 32542 482294
rect 31986 446378 32222 446614
rect 32306 446378 32542 446614
rect 31986 446058 32222 446294
rect 32306 446058 32542 446294
rect 31986 410378 32222 410614
rect 32306 410378 32542 410614
rect 31986 410058 32222 410294
rect 32306 410058 32542 410294
rect 31986 374378 32222 374614
rect 32306 374378 32542 374614
rect 31986 374058 32222 374294
rect 32306 374058 32542 374294
rect 31986 338378 32222 338614
rect 32306 338378 32542 338614
rect 31986 338058 32222 338294
rect 32306 338058 32542 338294
rect 31986 302378 32222 302614
rect 32306 302378 32542 302614
rect 31986 302058 32222 302294
rect 32306 302058 32542 302294
rect 31986 266378 32222 266614
rect 32306 266378 32542 266614
rect 31986 266058 32222 266294
rect 32306 266058 32542 266294
rect 31986 230378 32222 230614
rect 32306 230378 32542 230614
rect 31986 230058 32222 230294
rect 32306 230058 32542 230294
rect 31986 194378 32222 194614
rect 32306 194378 32542 194614
rect 31986 194058 32222 194294
rect 32306 194058 32542 194294
rect 31986 158378 32222 158614
rect 32306 158378 32542 158614
rect 31986 158058 32222 158294
rect 32306 158058 32542 158294
rect 31986 122378 32222 122614
rect 32306 122378 32542 122614
rect 31986 122058 32222 122294
rect 32306 122058 32542 122294
rect 31986 86378 32222 86614
rect 32306 86378 32542 86614
rect 31986 86058 32222 86294
rect 32306 86058 32542 86294
rect 34546 707482 34782 707718
rect 34866 707482 35102 707718
rect 34546 707162 34782 707398
rect 34866 707162 35102 707398
rect 34546 672938 34782 673174
rect 34866 672938 35102 673174
rect 34546 672618 34782 672854
rect 34866 672618 35102 672854
rect 34546 636938 34782 637174
rect 34866 636938 35102 637174
rect 34546 636618 34782 636854
rect 34866 636618 35102 636854
rect 34546 600938 34782 601174
rect 34866 600938 35102 601174
rect 34546 600618 34782 600854
rect 34866 600618 35102 600854
rect 34546 564938 34782 565174
rect 34866 564938 35102 565174
rect 34546 564618 34782 564854
rect 34866 564618 35102 564854
rect 34546 528938 34782 529174
rect 34866 528938 35102 529174
rect 34546 528618 34782 528854
rect 34866 528618 35102 528854
rect 34546 492938 34782 493174
rect 34866 492938 35102 493174
rect 34546 492618 34782 492854
rect 34866 492618 35102 492854
rect 34546 456938 34782 457174
rect 34866 456938 35102 457174
rect 34546 456618 34782 456854
rect 34866 456618 35102 456854
rect 34546 420938 34782 421174
rect 34866 420938 35102 421174
rect 34546 420618 34782 420854
rect 34866 420618 35102 420854
rect 34546 384938 34782 385174
rect 34866 384938 35102 385174
rect 34546 384618 34782 384854
rect 34866 384618 35102 384854
rect 34546 348938 34782 349174
rect 34866 348938 35102 349174
rect 34546 348618 34782 348854
rect 34866 348618 35102 348854
rect 34546 312938 34782 313174
rect 34866 312938 35102 313174
rect 34546 312618 34782 312854
rect 34866 312618 35102 312854
rect 34546 276938 34782 277174
rect 34866 276938 35102 277174
rect 34546 276618 34782 276854
rect 34866 276618 35102 276854
rect 34546 240938 34782 241174
rect 34866 240938 35102 241174
rect 34546 240618 34782 240854
rect 34866 240618 35102 240854
rect 34546 204938 34782 205174
rect 34866 204938 35102 205174
rect 34546 204618 34782 204854
rect 34866 204618 35102 204854
rect 34546 168938 34782 169174
rect 34866 168938 35102 169174
rect 34546 168618 34782 168854
rect 34866 168618 35102 168854
rect 34546 132938 34782 133174
rect 34866 132938 35102 133174
rect 34546 132618 34782 132854
rect 34866 132618 35102 132854
rect 34546 96938 34782 97174
rect 34866 96938 35102 97174
rect 34546 96618 34782 96854
rect 34866 96618 35102 96854
rect 38266 676658 38502 676894
rect 38586 676658 38822 676894
rect 38266 676338 38502 676574
rect 38586 676338 38822 676574
rect 38266 640658 38502 640894
rect 38586 640658 38822 640894
rect 38266 640338 38502 640574
rect 38586 640338 38822 640574
rect 38266 604658 38502 604894
rect 38586 604658 38822 604894
rect 38266 604338 38502 604574
rect 38586 604338 38822 604574
rect 38266 568658 38502 568894
rect 38586 568658 38822 568894
rect 38266 568338 38502 568574
rect 38586 568338 38822 568574
rect 38266 532658 38502 532894
rect 38586 532658 38822 532894
rect 38266 532338 38502 532574
rect 38586 532338 38822 532574
rect 38266 496658 38502 496894
rect 38586 496658 38822 496894
rect 38266 496338 38502 496574
rect 38586 496338 38822 496574
rect 38266 460658 38502 460894
rect 38586 460658 38822 460894
rect 38266 460338 38502 460574
rect 38586 460338 38822 460574
rect 38266 424658 38502 424894
rect 38586 424658 38822 424894
rect 38266 424338 38502 424574
rect 38586 424338 38822 424574
rect 38266 388658 38502 388894
rect 38586 388658 38822 388894
rect 38266 388338 38502 388574
rect 38586 388338 38822 388574
rect 38266 352658 38502 352894
rect 38586 352658 38822 352894
rect 38266 352338 38502 352574
rect 38586 352338 38822 352574
rect 38266 316658 38502 316894
rect 38586 316658 38822 316894
rect 38266 316338 38502 316574
rect 38586 316338 38822 316574
rect 38266 280658 38502 280894
rect 38586 280658 38822 280894
rect 38266 280338 38502 280574
rect 38586 280338 38822 280574
rect 38266 244658 38502 244894
rect 38586 244658 38822 244894
rect 38266 244338 38502 244574
rect 38586 244338 38822 244574
rect 38266 208658 38502 208894
rect 38586 208658 38822 208894
rect 38266 208338 38502 208574
rect 38586 208338 38822 208574
rect 38266 172658 38502 172894
rect 38586 172658 38822 172894
rect 38266 172338 38502 172574
rect 38586 172338 38822 172574
rect 38266 136658 38502 136894
rect 38586 136658 38822 136894
rect 38266 136338 38502 136574
rect 38586 136338 38822 136574
rect 38266 100658 38502 100894
rect 38586 100658 38822 100894
rect 38266 100338 38502 100574
rect 38586 100338 38822 100574
rect 40826 704602 41062 704838
rect 41146 704602 41382 704838
rect 40826 704282 41062 704518
rect 41146 704282 41382 704518
rect 40826 687218 41062 687454
rect 41146 687218 41382 687454
rect 40826 686898 41062 687134
rect 41146 686898 41382 687134
rect 40826 651218 41062 651454
rect 41146 651218 41382 651454
rect 40826 650898 41062 651134
rect 41146 650898 41382 651134
rect 40826 615218 41062 615454
rect 41146 615218 41382 615454
rect 40826 614898 41062 615134
rect 41146 614898 41382 615134
rect 40826 579218 41062 579454
rect 41146 579218 41382 579454
rect 40826 578898 41062 579134
rect 41146 578898 41382 579134
rect 40826 543218 41062 543454
rect 41146 543218 41382 543454
rect 40826 542898 41062 543134
rect 41146 542898 41382 543134
rect 40826 507218 41062 507454
rect 41146 507218 41382 507454
rect 40826 506898 41062 507134
rect 41146 506898 41382 507134
rect 40826 471218 41062 471454
rect 41146 471218 41382 471454
rect 40826 470898 41062 471134
rect 41146 470898 41382 471134
rect 40826 435218 41062 435454
rect 41146 435218 41382 435454
rect 40826 434898 41062 435134
rect 41146 434898 41382 435134
rect 40826 399218 41062 399454
rect 41146 399218 41382 399454
rect 40826 398898 41062 399134
rect 41146 398898 41382 399134
rect 40826 363218 41062 363454
rect 41146 363218 41382 363454
rect 40826 362898 41062 363134
rect 41146 362898 41382 363134
rect 40826 327218 41062 327454
rect 41146 327218 41382 327454
rect 40826 326898 41062 327134
rect 41146 326898 41382 327134
rect 40826 291218 41062 291454
rect 41146 291218 41382 291454
rect 40826 290898 41062 291134
rect 41146 290898 41382 291134
rect 40826 255218 41062 255454
rect 41146 255218 41382 255454
rect 40826 254898 41062 255134
rect 41146 254898 41382 255134
rect 40826 219218 41062 219454
rect 41146 219218 41382 219454
rect 40826 218898 41062 219134
rect 41146 218898 41382 219134
rect 40826 183218 41062 183454
rect 41146 183218 41382 183454
rect 40826 182898 41062 183134
rect 41146 182898 41382 183134
rect 40826 147218 41062 147454
rect 41146 147218 41382 147454
rect 40826 146898 41062 147134
rect 41146 146898 41382 147134
rect 40826 111218 41062 111454
rect 41146 111218 41382 111454
rect 40826 110898 41062 111134
rect 41146 110898 41382 111134
rect 40826 75218 41062 75454
rect 41146 75218 41382 75454
rect 40826 74898 41062 75134
rect 41146 74898 41382 75134
rect 51986 710362 52222 710598
rect 52306 710362 52542 710598
rect 51986 710042 52222 710278
rect 52306 710042 52542 710278
rect 48266 708442 48502 708678
rect 48586 708442 48822 708678
rect 48266 708122 48502 708358
rect 48586 708122 48822 708358
rect 41986 680378 42222 680614
rect 42306 680378 42542 680614
rect 41986 680058 42222 680294
rect 42306 680058 42542 680294
rect 41986 644378 42222 644614
rect 42306 644378 42542 644614
rect 41986 644058 42222 644294
rect 42306 644058 42542 644294
rect 41986 608378 42222 608614
rect 42306 608378 42542 608614
rect 41986 608058 42222 608294
rect 42306 608058 42542 608294
rect 41986 572378 42222 572614
rect 42306 572378 42542 572614
rect 41986 572058 42222 572294
rect 42306 572058 42542 572294
rect 41986 536378 42222 536614
rect 42306 536378 42542 536614
rect 41986 536058 42222 536294
rect 42306 536058 42542 536294
rect 41986 500378 42222 500614
rect 42306 500378 42542 500614
rect 41986 500058 42222 500294
rect 42306 500058 42542 500294
rect 41986 464378 42222 464614
rect 42306 464378 42542 464614
rect 41986 464058 42222 464294
rect 42306 464058 42542 464294
rect 41986 428378 42222 428614
rect 42306 428378 42542 428614
rect 41986 428058 42222 428294
rect 42306 428058 42542 428294
rect 41986 392378 42222 392614
rect 42306 392378 42542 392614
rect 41986 392058 42222 392294
rect 42306 392058 42542 392294
rect 41986 356378 42222 356614
rect 42306 356378 42542 356614
rect 41986 356058 42222 356294
rect 42306 356058 42542 356294
rect 41986 320378 42222 320614
rect 42306 320378 42542 320614
rect 41986 320058 42222 320294
rect 42306 320058 42542 320294
rect 41986 284378 42222 284614
rect 42306 284378 42542 284614
rect 41986 284058 42222 284294
rect 42306 284058 42542 284294
rect 41986 248378 42222 248614
rect 42306 248378 42542 248614
rect 41986 248058 42222 248294
rect 42306 248058 42542 248294
rect 41986 212378 42222 212614
rect 42306 212378 42542 212614
rect 41986 212058 42222 212294
rect 42306 212058 42542 212294
rect 41986 176378 42222 176614
rect 42306 176378 42542 176614
rect 41986 176058 42222 176294
rect 42306 176058 42542 176294
rect 41986 140378 42222 140614
rect 42306 140378 42542 140614
rect 41986 140058 42222 140294
rect 42306 140058 42542 140294
rect 41986 104378 42222 104614
rect 42306 104378 42542 104614
rect 41986 104058 42222 104294
rect 42306 104058 42542 104294
rect 44546 706522 44782 706758
rect 44866 706522 45102 706758
rect 44546 706202 44782 706438
rect 44866 706202 45102 706438
rect 44546 690938 44782 691174
rect 44866 690938 45102 691174
rect 44546 690618 44782 690854
rect 44866 690618 45102 690854
rect 44546 654938 44782 655174
rect 44866 654938 45102 655174
rect 44546 654618 44782 654854
rect 44866 654618 45102 654854
rect 44546 618938 44782 619174
rect 44866 618938 45102 619174
rect 44546 618618 44782 618854
rect 44866 618618 45102 618854
rect 44546 582938 44782 583174
rect 44866 582938 45102 583174
rect 44546 582618 44782 582854
rect 44866 582618 45102 582854
rect 44546 546938 44782 547174
rect 44866 546938 45102 547174
rect 44546 546618 44782 546854
rect 44866 546618 45102 546854
rect 44546 510938 44782 511174
rect 44866 510938 45102 511174
rect 44546 510618 44782 510854
rect 44866 510618 45102 510854
rect 44546 474938 44782 475174
rect 44866 474938 45102 475174
rect 44546 474618 44782 474854
rect 44866 474618 45102 474854
rect 44546 438938 44782 439174
rect 44866 438938 45102 439174
rect 44546 438618 44782 438854
rect 44866 438618 45102 438854
rect 44546 402938 44782 403174
rect 44866 402938 45102 403174
rect 44546 402618 44782 402854
rect 44866 402618 45102 402854
rect 44546 366938 44782 367174
rect 44866 366938 45102 367174
rect 44546 366618 44782 366854
rect 44866 366618 45102 366854
rect 44546 330938 44782 331174
rect 44866 330938 45102 331174
rect 44546 330618 44782 330854
rect 44866 330618 45102 330854
rect 44546 294938 44782 295174
rect 44866 294938 45102 295174
rect 44546 294618 44782 294854
rect 44866 294618 45102 294854
rect 44546 258938 44782 259174
rect 44866 258938 45102 259174
rect 44546 258618 44782 258854
rect 44866 258618 45102 258854
rect 44546 222938 44782 223174
rect 44866 222938 45102 223174
rect 44546 222618 44782 222854
rect 44866 222618 45102 222854
rect 44546 186938 44782 187174
rect 44866 186938 45102 187174
rect 44546 186618 44782 186854
rect 44866 186618 45102 186854
rect 44546 150938 44782 151174
rect 44866 150938 45102 151174
rect 44546 150618 44782 150854
rect 44866 150618 45102 150854
rect 44546 114938 44782 115174
rect 44866 114938 45102 115174
rect 44546 114618 44782 114854
rect 44866 114618 45102 114854
rect 44546 78938 44782 79174
rect 44866 78938 45102 79174
rect 44546 78618 44782 78854
rect 44866 78618 45102 78854
rect 48266 694658 48502 694894
rect 48586 694658 48822 694894
rect 48266 694338 48502 694574
rect 48586 694338 48822 694574
rect 48266 658658 48502 658894
rect 48586 658658 48822 658894
rect 48266 658338 48502 658574
rect 48586 658338 48822 658574
rect 48266 622658 48502 622894
rect 48586 622658 48822 622894
rect 48266 622338 48502 622574
rect 48586 622338 48822 622574
rect 48266 586658 48502 586894
rect 48586 586658 48822 586894
rect 48266 586338 48502 586574
rect 48586 586338 48822 586574
rect 48266 550658 48502 550894
rect 48586 550658 48822 550894
rect 48266 550338 48502 550574
rect 48586 550338 48822 550574
rect 48266 514658 48502 514894
rect 48586 514658 48822 514894
rect 48266 514338 48502 514574
rect 48586 514338 48822 514574
rect 48266 478658 48502 478894
rect 48586 478658 48822 478894
rect 48266 478338 48502 478574
rect 48586 478338 48822 478574
rect 48266 442658 48502 442894
rect 48586 442658 48822 442894
rect 48266 442338 48502 442574
rect 48586 442338 48822 442574
rect 48266 406658 48502 406894
rect 48586 406658 48822 406894
rect 48266 406338 48502 406574
rect 48586 406338 48822 406574
rect 48266 370658 48502 370894
rect 48586 370658 48822 370894
rect 48266 370338 48502 370574
rect 48586 370338 48822 370574
rect 48266 334658 48502 334894
rect 48586 334658 48822 334894
rect 48266 334338 48502 334574
rect 48586 334338 48822 334574
rect 48266 298658 48502 298894
rect 48586 298658 48822 298894
rect 48266 298338 48502 298574
rect 48586 298338 48822 298574
rect 48266 262658 48502 262894
rect 48586 262658 48822 262894
rect 48266 262338 48502 262574
rect 48586 262338 48822 262574
rect 48266 226658 48502 226894
rect 48586 226658 48822 226894
rect 48266 226338 48502 226574
rect 48586 226338 48822 226574
rect 48266 190658 48502 190894
rect 48586 190658 48822 190894
rect 48266 190338 48502 190574
rect 48586 190338 48822 190574
rect 48266 154658 48502 154894
rect 48586 154658 48822 154894
rect 48266 154338 48502 154574
rect 48586 154338 48822 154574
rect 48266 118658 48502 118894
rect 48586 118658 48822 118894
rect 48266 118338 48502 118574
rect 48586 118338 48822 118574
rect 48266 82658 48502 82894
rect 48586 82658 48822 82894
rect 48266 82338 48502 82574
rect 48586 82338 48822 82574
rect 50826 705562 51062 705798
rect 51146 705562 51382 705798
rect 50826 705242 51062 705478
rect 51146 705242 51382 705478
rect 50826 669218 51062 669454
rect 51146 669218 51382 669454
rect 50826 668898 51062 669134
rect 51146 668898 51382 669134
rect 50826 633218 51062 633454
rect 51146 633218 51382 633454
rect 50826 632898 51062 633134
rect 51146 632898 51382 633134
rect 50826 597218 51062 597454
rect 51146 597218 51382 597454
rect 50826 596898 51062 597134
rect 51146 596898 51382 597134
rect 50826 561218 51062 561454
rect 51146 561218 51382 561454
rect 50826 560898 51062 561134
rect 51146 560898 51382 561134
rect 50826 525218 51062 525454
rect 51146 525218 51382 525454
rect 50826 524898 51062 525134
rect 51146 524898 51382 525134
rect 50826 489218 51062 489454
rect 51146 489218 51382 489454
rect 50826 488898 51062 489134
rect 51146 488898 51382 489134
rect 50826 453218 51062 453454
rect 51146 453218 51382 453454
rect 50826 452898 51062 453134
rect 51146 452898 51382 453134
rect 50826 417218 51062 417454
rect 51146 417218 51382 417454
rect 50826 416898 51062 417134
rect 51146 416898 51382 417134
rect 50826 381218 51062 381454
rect 51146 381218 51382 381454
rect 50826 380898 51062 381134
rect 51146 380898 51382 381134
rect 50826 345218 51062 345454
rect 51146 345218 51382 345454
rect 50826 344898 51062 345134
rect 51146 344898 51382 345134
rect 50826 309218 51062 309454
rect 51146 309218 51382 309454
rect 50826 308898 51062 309134
rect 51146 308898 51382 309134
rect 50826 273218 51062 273454
rect 51146 273218 51382 273454
rect 50826 272898 51062 273134
rect 51146 272898 51382 273134
rect 50826 237218 51062 237454
rect 51146 237218 51382 237454
rect 50826 236898 51062 237134
rect 51146 236898 51382 237134
rect 50826 201218 51062 201454
rect 51146 201218 51382 201454
rect 50826 200898 51062 201134
rect 51146 200898 51382 201134
rect 50826 165218 51062 165454
rect 51146 165218 51382 165454
rect 50826 164898 51062 165134
rect 51146 164898 51382 165134
rect 50826 129218 51062 129454
rect 51146 129218 51382 129454
rect 50826 128898 51062 129134
rect 51146 128898 51382 129134
rect 50826 93218 51062 93454
rect 51146 93218 51382 93454
rect 50826 92898 51062 93134
rect 51146 92898 51382 93134
rect 61986 711322 62222 711558
rect 62306 711322 62542 711558
rect 61986 711002 62222 711238
rect 62306 711002 62542 711238
rect 58266 709402 58502 709638
rect 58586 709402 58822 709638
rect 58266 709082 58502 709318
rect 58586 709082 58822 709318
rect 51986 698378 52222 698614
rect 52306 698378 52542 698614
rect 51986 698058 52222 698294
rect 52306 698058 52542 698294
rect 51986 662378 52222 662614
rect 52306 662378 52542 662614
rect 51986 662058 52222 662294
rect 52306 662058 52542 662294
rect 51986 626378 52222 626614
rect 52306 626378 52542 626614
rect 51986 626058 52222 626294
rect 52306 626058 52542 626294
rect 51986 590378 52222 590614
rect 52306 590378 52542 590614
rect 51986 590058 52222 590294
rect 52306 590058 52542 590294
rect 51986 554378 52222 554614
rect 52306 554378 52542 554614
rect 51986 554058 52222 554294
rect 52306 554058 52542 554294
rect 51986 518378 52222 518614
rect 52306 518378 52542 518614
rect 51986 518058 52222 518294
rect 52306 518058 52542 518294
rect 51986 482378 52222 482614
rect 52306 482378 52542 482614
rect 51986 482058 52222 482294
rect 52306 482058 52542 482294
rect 51986 446378 52222 446614
rect 52306 446378 52542 446614
rect 51986 446058 52222 446294
rect 52306 446058 52542 446294
rect 51986 410378 52222 410614
rect 52306 410378 52542 410614
rect 51986 410058 52222 410294
rect 52306 410058 52542 410294
rect 51986 374378 52222 374614
rect 52306 374378 52542 374614
rect 51986 374058 52222 374294
rect 52306 374058 52542 374294
rect 51986 338378 52222 338614
rect 52306 338378 52542 338614
rect 51986 338058 52222 338294
rect 52306 338058 52542 338294
rect 51986 302378 52222 302614
rect 52306 302378 52542 302614
rect 51986 302058 52222 302294
rect 52306 302058 52542 302294
rect 51986 266378 52222 266614
rect 52306 266378 52542 266614
rect 51986 266058 52222 266294
rect 52306 266058 52542 266294
rect 51986 230378 52222 230614
rect 52306 230378 52542 230614
rect 51986 230058 52222 230294
rect 52306 230058 52542 230294
rect 51986 194378 52222 194614
rect 52306 194378 52542 194614
rect 51986 194058 52222 194294
rect 52306 194058 52542 194294
rect 51986 158378 52222 158614
rect 52306 158378 52542 158614
rect 51986 158058 52222 158294
rect 52306 158058 52542 158294
rect 51986 122378 52222 122614
rect 52306 122378 52542 122614
rect 51986 122058 52222 122294
rect 52306 122058 52542 122294
rect 51986 86378 52222 86614
rect 52306 86378 52542 86614
rect 51986 86058 52222 86294
rect 52306 86058 52542 86294
rect 54546 707482 54782 707718
rect 54866 707482 55102 707718
rect 54546 707162 54782 707398
rect 54866 707162 55102 707398
rect 54546 672938 54782 673174
rect 54866 672938 55102 673174
rect 54546 672618 54782 672854
rect 54866 672618 55102 672854
rect 54546 636938 54782 637174
rect 54866 636938 55102 637174
rect 54546 636618 54782 636854
rect 54866 636618 55102 636854
rect 54546 600938 54782 601174
rect 54866 600938 55102 601174
rect 54546 600618 54782 600854
rect 54866 600618 55102 600854
rect 54546 564938 54782 565174
rect 54866 564938 55102 565174
rect 54546 564618 54782 564854
rect 54866 564618 55102 564854
rect 54546 528938 54782 529174
rect 54866 528938 55102 529174
rect 54546 528618 54782 528854
rect 54866 528618 55102 528854
rect 54546 492938 54782 493174
rect 54866 492938 55102 493174
rect 54546 492618 54782 492854
rect 54866 492618 55102 492854
rect 54546 456938 54782 457174
rect 54866 456938 55102 457174
rect 54546 456618 54782 456854
rect 54866 456618 55102 456854
rect 54546 420938 54782 421174
rect 54866 420938 55102 421174
rect 54546 420618 54782 420854
rect 54866 420618 55102 420854
rect 54546 384938 54782 385174
rect 54866 384938 55102 385174
rect 54546 384618 54782 384854
rect 54866 384618 55102 384854
rect 54546 348938 54782 349174
rect 54866 348938 55102 349174
rect 54546 348618 54782 348854
rect 54866 348618 55102 348854
rect 54546 312938 54782 313174
rect 54866 312938 55102 313174
rect 54546 312618 54782 312854
rect 54866 312618 55102 312854
rect 54546 276938 54782 277174
rect 54866 276938 55102 277174
rect 54546 276618 54782 276854
rect 54866 276618 55102 276854
rect 54546 240938 54782 241174
rect 54866 240938 55102 241174
rect 54546 240618 54782 240854
rect 54866 240618 55102 240854
rect 54546 204938 54782 205174
rect 54866 204938 55102 205174
rect 54546 204618 54782 204854
rect 54866 204618 55102 204854
rect 54546 168938 54782 169174
rect 54866 168938 55102 169174
rect 54546 168618 54782 168854
rect 54866 168618 55102 168854
rect 54546 132938 54782 133174
rect 54866 132938 55102 133174
rect 54546 132618 54782 132854
rect 54866 132618 55102 132854
rect 54546 96938 54782 97174
rect 54866 96938 55102 97174
rect 54546 96618 54782 96854
rect 54866 96618 55102 96854
rect 58266 676658 58502 676894
rect 58586 676658 58822 676894
rect 58266 676338 58502 676574
rect 58586 676338 58822 676574
rect 58266 640658 58502 640894
rect 58586 640658 58822 640894
rect 58266 640338 58502 640574
rect 58586 640338 58822 640574
rect 58266 604658 58502 604894
rect 58586 604658 58822 604894
rect 58266 604338 58502 604574
rect 58586 604338 58822 604574
rect 58266 568658 58502 568894
rect 58586 568658 58822 568894
rect 58266 568338 58502 568574
rect 58586 568338 58822 568574
rect 58266 532658 58502 532894
rect 58586 532658 58822 532894
rect 58266 532338 58502 532574
rect 58586 532338 58822 532574
rect 58266 496658 58502 496894
rect 58586 496658 58822 496894
rect 58266 496338 58502 496574
rect 58586 496338 58822 496574
rect 58266 460658 58502 460894
rect 58586 460658 58822 460894
rect 58266 460338 58502 460574
rect 58586 460338 58822 460574
rect 58266 424658 58502 424894
rect 58586 424658 58822 424894
rect 58266 424338 58502 424574
rect 58586 424338 58822 424574
rect 58266 388658 58502 388894
rect 58586 388658 58822 388894
rect 58266 388338 58502 388574
rect 58586 388338 58822 388574
rect 58266 352658 58502 352894
rect 58586 352658 58822 352894
rect 58266 352338 58502 352574
rect 58586 352338 58822 352574
rect 58266 316658 58502 316894
rect 58586 316658 58822 316894
rect 58266 316338 58502 316574
rect 58586 316338 58822 316574
rect 58266 280658 58502 280894
rect 58586 280658 58822 280894
rect 58266 280338 58502 280574
rect 58586 280338 58822 280574
rect 58266 244658 58502 244894
rect 58586 244658 58822 244894
rect 58266 244338 58502 244574
rect 58586 244338 58822 244574
rect 58266 208658 58502 208894
rect 58586 208658 58822 208894
rect 58266 208338 58502 208574
rect 58586 208338 58822 208574
rect 58266 172658 58502 172894
rect 58586 172658 58822 172894
rect 58266 172338 58502 172574
rect 58586 172338 58822 172574
rect 58266 136658 58502 136894
rect 58586 136658 58822 136894
rect 58266 136338 58502 136574
rect 58586 136338 58822 136574
rect 58266 100658 58502 100894
rect 58586 100658 58822 100894
rect 58266 100338 58502 100574
rect 58586 100338 58822 100574
rect 60826 704602 61062 704838
rect 61146 704602 61382 704838
rect 60826 704282 61062 704518
rect 61146 704282 61382 704518
rect 60826 687218 61062 687454
rect 61146 687218 61382 687454
rect 60826 686898 61062 687134
rect 61146 686898 61382 687134
rect 60826 651218 61062 651454
rect 61146 651218 61382 651454
rect 60826 650898 61062 651134
rect 61146 650898 61382 651134
rect 60826 615218 61062 615454
rect 61146 615218 61382 615454
rect 60826 614898 61062 615134
rect 61146 614898 61382 615134
rect 60826 579218 61062 579454
rect 61146 579218 61382 579454
rect 60826 578898 61062 579134
rect 61146 578898 61382 579134
rect 60826 543218 61062 543454
rect 61146 543218 61382 543454
rect 60826 542898 61062 543134
rect 61146 542898 61382 543134
rect 60826 507218 61062 507454
rect 61146 507218 61382 507454
rect 60826 506898 61062 507134
rect 61146 506898 61382 507134
rect 60826 471218 61062 471454
rect 61146 471218 61382 471454
rect 60826 470898 61062 471134
rect 61146 470898 61382 471134
rect 60826 435218 61062 435454
rect 61146 435218 61382 435454
rect 60826 434898 61062 435134
rect 61146 434898 61382 435134
rect 60826 399218 61062 399454
rect 61146 399218 61382 399454
rect 60826 398898 61062 399134
rect 61146 398898 61382 399134
rect 60826 363218 61062 363454
rect 61146 363218 61382 363454
rect 60826 362898 61062 363134
rect 61146 362898 61382 363134
rect 60826 327218 61062 327454
rect 61146 327218 61382 327454
rect 60826 326898 61062 327134
rect 61146 326898 61382 327134
rect 60826 291218 61062 291454
rect 61146 291218 61382 291454
rect 60826 290898 61062 291134
rect 61146 290898 61382 291134
rect 60826 255218 61062 255454
rect 61146 255218 61382 255454
rect 60826 254898 61062 255134
rect 61146 254898 61382 255134
rect 60826 219218 61062 219454
rect 61146 219218 61382 219454
rect 60826 218898 61062 219134
rect 61146 218898 61382 219134
rect 60826 183218 61062 183454
rect 61146 183218 61382 183454
rect 60826 182898 61062 183134
rect 61146 182898 61382 183134
rect 60826 147218 61062 147454
rect 61146 147218 61382 147454
rect 60826 146898 61062 147134
rect 61146 146898 61382 147134
rect 60826 111218 61062 111454
rect 61146 111218 61382 111454
rect 60826 110898 61062 111134
rect 61146 110898 61382 111134
rect 60826 75218 61062 75454
rect 61146 75218 61382 75454
rect 60826 74898 61062 75134
rect 61146 74898 61382 75134
rect 71986 710362 72222 710598
rect 72306 710362 72542 710598
rect 71986 710042 72222 710278
rect 72306 710042 72542 710278
rect 68266 708442 68502 708678
rect 68586 708442 68822 708678
rect 68266 708122 68502 708358
rect 68586 708122 68822 708358
rect 61986 680378 62222 680614
rect 62306 680378 62542 680614
rect 61986 680058 62222 680294
rect 62306 680058 62542 680294
rect 61986 644378 62222 644614
rect 62306 644378 62542 644614
rect 61986 644058 62222 644294
rect 62306 644058 62542 644294
rect 61986 608378 62222 608614
rect 62306 608378 62542 608614
rect 61986 608058 62222 608294
rect 62306 608058 62542 608294
rect 61986 572378 62222 572614
rect 62306 572378 62542 572614
rect 61986 572058 62222 572294
rect 62306 572058 62542 572294
rect 61986 536378 62222 536614
rect 62306 536378 62542 536614
rect 61986 536058 62222 536294
rect 62306 536058 62542 536294
rect 61986 500378 62222 500614
rect 62306 500378 62542 500614
rect 61986 500058 62222 500294
rect 62306 500058 62542 500294
rect 61986 464378 62222 464614
rect 62306 464378 62542 464614
rect 61986 464058 62222 464294
rect 62306 464058 62542 464294
rect 61986 428378 62222 428614
rect 62306 428378 62542 428614
rect 61986 428058 62222 428294
rect 62306 428058 62542 428294
rect 61986 392378 62222 392614
rect 62306 392378 62542 392614
rect 61986 392058 62222 392294
rect 62306 392058 62542 392294
rect 61986 356378 62222 356614
rect 62306 356378 62542 356614
rect 61986 356058 62222 356294
rect 62306 356058 62542 356294
rect 61986 320378 62222 320614
rect 62306 320378 62542 320614
rect 61986 320058 62222 320294
rect 62306 320058 62542 320294
rect 61986 284378 62222 284614
rect 62306 284378 62542 284614
rect 61986 284058 62222 284294
rect 62306 284058 62542 284294
rect 61986 248378 62222 248614
rect 62306 248378 62542 248614
rect 61986 248058 62222 248294
rect 62306 248058 62542 248294
rect 61986 212378 62222 212614
rect 62306 212378 62542 212614
rect 61986 212058 62222 212294
rect 62306 212058 62542 212294
rect 61986 176378 62222 176614
rect 62306 176378 62542 176614
rect 61986 176058 62222 176294
rect 62306 176058 62542 176294
rect 61986 140378 62222 140614
rect 62306 140378 62542 140614
rect 61986 140058 62222 140294
rect 62306 140058 62542 140294
rect 61986 104378 62222 104614
rect 62306 104378 62542 104614
rect 61986 104058 62222 104294
rect 62306 104058 62542 104294
rect 64546 706522 64782 706758
rect 64866 706522 65102 706758
rect 64546 706202 64782 706438
rect 64866 706202 65102 706438
rect 64546 690938 64782 691174
rect 64866 690938 65102 691174
rect 64546 690618 64782 690854
rect 64866 690618 65102 690854
rect 64546 654938 64782 655174
rect 64866 654938 65102 655174
rect 64546 654618 64782 654854
rect 64866 654618 65102 654854
rect 64546 618938 64782 619174
rect 64866 618938 65102 619174
rect 64546 618618 64782 618854
rect 64866 618618 65102 618854
rect 64546 582938 64782 583174
rect 64866 582938 65102 583174
rect 64546 582618 64782 582854
rect 64866 582618 65102 582854
rect 64546 546938 64782 547174
rect 64866 546938 65102 547174
rect 64546 546618 64782 546854
rect 64866 546618 65102 546854
rect 64546 510938 64782 511174
rect 64866 510938 65102 511174
rect 64546 510618 64782 510854
rect 64866 510618 65102 510854
rect 64546 474938 64782 475174
rect 64866 474938 65102 475174
rect 64546 474618 64782 474854
rect 64866 474618 65102 474854
rect 64546 438938 64782 439174
rect 64866 438938 65102 439174
rect 64546 438618 64782 438854
rect 64866 438618 65102 438854
rect 64546 402938 64782 403174
rect 64866 402938 65102 403174
rect 64546 402618 64782 402854
rect 64866 402618 65102 402854
rect 64546 366938 64782 367174
rect 64866 366938 65102 367174
rect 64546 366618 64782 366854
rect 64866 366618 65102 366854
rect 64546 330938 64782 331174
rect 64866 330938 65102 331174
rect 64546 330618 64782 330854
rect 64866 330618 65102 330854
rect 64546 294938 64782 295174
rect 64866 294938 65102 295174
rect 64546 294618 64782 294854
rect 64866 294618 65102 294854
rect 64546 258938 64782 259174
rect 64866 258938 65102 259174
rect 64546 258618 64782 258854
rect 64866 258618 65102 258854
rect 64546 222938 64782 223174
rect 64866 222938 65102 223174
rect 64546 222618 64782 222854
rect 64866 222618 65102 222854
rect 64546 186938 64782 187174
rect 64866 186938 65102 187174
rect 64546 186618 64782 186854
rect 64866 186618 65102 186854
rect 64546 150938 64782 151174
rect 64866 150938 65102 151174
rect 64546 150618 64782 150854
rect 64866 150618 65102 150854
rect 64546 114938 64782 115174
rect 64866 114938 65102 115174
rect 64546 114618 64782 114854
rect 64866 114618 65102 114854
rect 64546 78938 64782 79174
rect 64866 78938 65102 79174
rect 64546 78618 64782 78854
rect 64866 78618 65102 78854
rect 68266 694658 68502 694894
rect 68586 694658 68822 694894
rect 68266 694338 68502 694574
rect 68586 694338 68822 694574
rect 68266 658658 68502 658894
rect 68586 658658 68822 658894
rect 68266 658338 68502 658574
rect 68586 658338 68822 658574
rect 68266 622658 68502 622894
rect 68586 622658 68822 622894
rect 68266 622338 68502 622574
rect 68586 622338 68822 622574
rect 68266 586658 68502 586894
rect 68586 586658 68822 586894
rect 68266 586338 68502 586574
rect 68586 586338 68822 586574
rect 68266 550658 68502 550894
rect 68586 550658 68822 550894
rect 68266 550338 68502 550574
rect 68586 550338 68822 550574
rect 68266 514658 68502 514894
rect 68586 514658 68822 514894
rect 68266 514338 68502 514574
rect 68586 514338 68822 514574
rect 68266 478658 68502 478894
rect 68586 478658 68822 478894
rect 68266 478338 68502 478574
rect 68586 478338 68822 478574
rect 68266 442658 68502 442894
rect 68586 442658 68822 442894
rect 68266 442338 68502 442574
rect 68586 442338 68822 442574
rect 68266 406658 68502 406894
rect 68586 406658 68822 406894
rect 68266 406338 68502 406574
rect 68586 406338 68822 406574
rect 68266 370658 68502 370894
rect 68586 370658 68822 370894
rect 68266 370338 68502 370574
rect 68586 370338 68822 370574
rect 68266 334658 68502 334894
rect 68586 334658 68822 334894
rect 68266 334338 68502 334574
rect 68586 334338 68822 334574
rect 68266 298658 68502 298894
rect 68586 298658 68822 298894
rect 68266 298338 68502 298574
rect 68586 298338 68822 298574
rect 68266 262658 68502 262894
rect 68586 262658 68822 262894
rect 68266 262338 68502 262574
rect 68586 262338 68822 262574
rect 68266 226658 68502 226894
rect 68586 226658 68822 226894
rect 68266 226338 68502 226574
rect 68586 226338 68822 226574
rect 68266 190658 68502 190894
rect 68586 190658 68822 190894
rect 68266 190338 68502 190574
rect 68586 190338 68822 190574
rect 68266 154658 68502 154894
rect 68586 154658 68822 154894
rect 68266 154338 68502 154574
rect 68586 154338 68822 154574
rect 68266 118658 68502 118894
rect 68586 118658 68822 118894
rect 68266 118338 68502 118574
rect 68586 118338 68822 118574
rect 68266 82658 68502 82894
rect 68586 82658 68822 82894
rect 68266 82338 68502 82574
rect 68586 82338 68822 82574
rect 70826 705562 71062 705798
rect 71146 705562 71382 705798
rect 70826 705242 71062 705478
rect 71146 705242 71382 705478
rect 70826 669218 71062 669454
rect 71146 669218 71382 669454
rect 70826 668898 71062 669134
rect 71146 668898 71382 669134
rect 70826 633218 71062 633454
rect 71146 633218 71382 633454
rect 70826 632898 71062 633134
rect 71146 632898 71382 633134
rect 70826 597218 71062 597454
rect 71146 597218 71382 597454
rect 70826 596898 71062 597134
rect 71146 596898 71382 597134
rect 70826 561218 71062 561454
rect 71146 561218 71382 561454
rect 70826 560898 71062 561134
rect 71146 560898 71382 561134
rect 70826 525218 71062 525454
rect 71146 525218 71382 525454
rect 70826 524898 71062 525134
rect 71146 524898 71382 525134
rect 70826 489218 71062 489454
rect 71146 489218 71382 489454
rect 70826 488898 71062 489134
rect 71146 488898 71382 489134
rect 70826 453218 71062 453454
rect 71146 453218 71382 453454
rect 70826 452898 71062 453134
rect 71146 452898 71382 453134
rect 70826 417218 71062 417454
rect 71146 417218 71382 417454
rect 70826 416898 71062 417134
rect 71146 416898 71382 417134
rect 70826 381218 71062 381454
rect 71146 381218 71382 381454
rect 70826 380898 71062 381134
rect 71146 380898 71382 381134
rect 70826 345218 71062 345454
rect 71146 345218 71382 345454
rect 70826 344898 71062 345134
rect 71146 344898 71382 345134
rect 70826 309218 71062 309454
rect 71146 309218 71382 309454
rect 70826 308898 71062 309134
rect 71146 308898 71382 309134
rect 70826 273218 71062 273454
rect 71146 273218 71382 273454
rect 70826 272898 71062 273134
rect 71146 272898 71382 273134
rect 70826 237218 71062 237454
rect 71146 237218 71382 237454
rect 70826 236898 71062 237134
rect 71146 236898 71382 237134
rect 70826 201218 71062 201454
rect 71146 201218 71382 201454
rect 70826 200898 71062 201134
rect 71146 200898 71382 201134
rect 70826 165218 71062 165454
rect 71146 165218 71382 165454
rect 70826 164898 71062 165134
rect 71146 164898 71382 165134
rect 70826 129218 71062 129454
rect 71146 129218 71382 129454
rect 70826 128898 71062 129134
rect 71146 128898 71382 129134
rect 70826 93218 71062 93454
rect 71146 93218 71382 93454
rect 70826 92898 71062 93134
rect 71146 92898 71382 93134
rect 81986 711322 82222 711558
rect 82306 711322 82542 711558
rect 81986 711002 82222 711238
rect 82306 711002 82542 711238
rect 78266 709402 78502 709638
rect 78586 709402 78822 709638
rect 78266 709082 78502 709318
rect 78586 709082 78822 709318
rect 71986 698378 72222 698614
rect 72306 698378 72542 698614
rect 71986 698058 72222 698294
rect 72306 698058 72542 698294
rect 71986 662378 72222 662614
rect 72306 662378 72542 662614
rect 71986 662058 72222 662294
rect 72306 662058 72542 662294
rect 71986 626378 72222 626614
rect 72306 626378 72542 626614
rect 71986 626058 72222 626294
rect 72306 626058 72542 626294
rect 71986 590378 72222 590614
rect 72306 590378 72542 590614
rect 71986 590058 72222 590294
rect 72306 590058 72542 590294
rect 71986 554378 72222 554614
rect 72306 554378 72542 554614
rect 71986 554058 72222 554294
rect 72306 554058 72542 554294
rect 71986 518378 72222 518614
rect 72306 518378 72542 518614
rect 71986 518058 72222 518294
rect 72306 518058 72542 518294
rect 71986 482378 72222 482614
rect 72306 482378 72542 482614
rect 71986 482058 72222 482294
rect 72306 482058 72542 482294
rect 71986 446378 72222 446614
rect 72306 446378 72542 446614
rect 71986 446058 72222 446294
rect 72306 446058 72542 446294
rect 71986 410378 72222 410614
rect 72306 410378 72542 410614
rect 71986 410058 72222 410294
rect 72306 410058 72542 410294
rect 71986 374378 72222 374614
rect 72306 374378 72542 374614
rect 71986 374058 72222 374294
rect 72306 374058 72542 374294
rect 71986 338378 72222 338614
rect 72306 338378 72542 338614
rect 71986 338058 72222 338294
rect 72306 338058 72542 338294
rect 71986 302378 72222 302614
rect 72306 302378 72542 302614
rect 71986 302058 72222 302294
rect 72306 302058 72542 302294
rect 71986 266378 72222 266614
rect 72306 266378 72542 266614
rect 71986 266058 72222 266294
rect 72306 266058 72542 266294
rect 71986 230378 72222 230614
rect 72306 230378 72542 230614
rect 71986 230058 72222 230294
rect 72306 230058 72542 230294
rect 71986 194378 72222 194614
rect 72306 194378 72542 194614
rect 71986 194058 72222 194294
rect 72306 194058 72542 194294
rect 71986 158378 72222 158614
rect 72306 158378 72542 158614
rect 71986 158058 72222 158294
rect 72306 158058 72542 158294
rect 71986 122378 72222 122614
rect 72306 122378 72542 122614
rect 71986 122058 72222 122294
rect 72306 122058 72542 122294
rect 71986 86378 72222 86614
rect 72306 86378 72542 86614
rect 71986 86058 72222 86294
rect 72306 86058 72542 86294
rect 74546 707482 74782 707718
rect 74866 707482 75102 707718
rect 74546 707162 74782 707398
rect 74866 707162 75102 707398
rect 74546 672938 74782 673174
rect 74866 672938 75102 673174
rect 74546 672618 74782 672854
rect 74866 672618 75102 672854
rect 74546 636938 74782 637174
rect 74866 636938 75102 637174
rect 74546 636618 74782 636854
rect 74866 636618 75102 636854
rect 74546 600938 74782 601174
rect 74866 600938 75102 601174
rect 74546 600618 74782 600854
rect 74866 600618 75102 600854
rect 74546 564938 74782 565174
rect 74866 564938 75102 565174
rect 74546 564618 74782 564854
rect 74866 564618 75102 564854
rect 74546 528938 74782 529174
rect 74866 528938 75102 529174
rect 74546 528618 74782 528854
rect 74866 528618 75102 528854
rect 74546 492938 74782 493174
rect 74866 492938 75102 493174
rect 74546 492618 74782 492854
rect 74866 492618 75102 492854
rect 74546 456938 74782 457174
rect 74866 456938 75102 457174
rect 74546 456618 74782 456854
rect 74866 456618 75102 456854
rect 74546 420938 74782 421174
rect 74866 420938 75102 421174
rect 74546 420618 74782 420854
rect 74866 420618 75102 420854
rect 74546 384938 74782 385174
rect 74866 384938 75102 385174
rect 74546 384618 74782 384854
rect 74866 384618 75102 384854
rect 74546 348938 74782 349174
rect 74866 348938 75102 349174
rect 74546 348618 74782 348854
rect 74866 348618 75102 348854
rect 74546 312938 74782 313174
rect 74866 312938 75102 313174
rect 74546 312618 74782 312854
rect 74866 312618 75102 312854
rect 74546 276938 74782 277174
rect 74866 276938 75102 277174
rect 74546 276618 74782 276854
rect 74866 276618 75102 276854
rect 74546 240938 74782 241174
rect 74866 240938 75102 241174
rect 74546 240618 74782 240854
rect 74866 240618 75102 240854
rect 74546 204938 74782 205174
rect 74866 204938 75102 205174
rect 74546 204618 74782 204854
rect 74866 204618 75102 204854
rect 74546 168938 74782 169174
rect 74866 168938 75102 169174
rect 74546 168618 74782 168854
rect 74866 168618 75102 168854
rect 74546 132938 74782 133174
rect 74866 132938 75102 133174
rect 74546 132618 74782 132854
rect 74866 132618 75102 132854
rect 74546 96938 74782 97174
rect 74866 96938 75102 97174
rect 74546 96618 74782 96854
rect 74866 96618 75102 96854
rect 14546 60938 14782 61174
rect 14866 60938 15102 61174
rect 14546 60618 14782 60854
rect 14866 60618 15102 60854
rect 24250 39218 24486 39454
rect 24250 38898 24486 39134
rect 14546 24938 14782 25174
rect 14866 24938 15102 25174
rect 14546 24618 14782 24854
rect 14866 24618 15102 24854
rect 14546 -3462 14782 -3226
rect 14866 -3462 15102 -3226
rect 14546 -3782 14782 -3546
rect 14866 -3782 15102 -3546
rect 20826 3218 21062 3454
rect 21146 3218 21382 3454
rect 20826 2898 21062 3134
rect 21146 2898 21382 3134
rect 20826 -582 21062 -346
rect 21146 -582 21382 -346
rect 20826 -902 21062 -666
rect 21146 -902 21382 -666
rect 18266 -5382 18502 -5146
rect 18586 -5382 18822 -5146
rect 18266 -5702 18502 -5466
rect 18586 -5702 18822 -5466
rect 11986 -6342 12222 -6106
rect 12306 -6342 12542 -6106
rect 11986 -6662 12222 -6426
rect 12306 -6662 12542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 24546 6938 24782 7174
rect 24866 6938 25102 7174
rect 24546 6618 24782 6854
rect 24866 6618 25102 6854
rect 24546 -2502 24782 -2266
rect 24866 -2502 25102 -2266
rect 24546 -2822 24782 -2586
rect 24866 -2822 25102 -2586
rect 28266 10658 28502 10894
rect 28586 10658 28822 10894
rect 28266 10338 28502 10574
rect 28586 10338 28822 10574
rect 74546 60938 74782 61174
rect 74866 60938 75102 61174
rect 74546 60618 74782 60854
rect 74866 60618 75102 60854
rect 39610 57218 39846 57454
rect 39610 56898 39846 57134
rect 54970 39218 55206 39454
rect 54970 38898 55206 39134
rect 74546 24938 74782 25174
rect 74866 24938 75102 25174
rect 74546 24618 74782 24854
rect 74866 24618 75102 24854
rect 31986 14378 32222 14614
rect 32306 14378 32542 14614
rect 31986 14058 32222 14294
rect 32306 14058 32542 14294
rect 30826 -1542 31062 -1306
rect 31146 -1542 31382 -1306
rect 30826 -1862 31062 -1626
rect 31146 -1862 31382 -1626
rect 28266 -4422 28502 -4186
rect 28586 -4422 28822 -4186
rect 28266 -4742 28502 -4506
rect 28586 -4742 28822 -4506
rect 21986 -7302 22222 -7066
rect 22306 -7302 22542 -7066
rect 21986 -7622 22222 -7386
rect 22306 -7622 22542 -7386
rect 34546 -3462 34782 -3226
rect 34866 -3462 35102 -3226
rect 34546 -3782 34782 -3546
rect 34866 -3782 35102 -3546
rect 40826 3218 41062 3454
rect 41146 3218 41382 3454
rect 40826 2898 41062 3134
rect 41146 2898 41382 3134
rect 40826 -582 41062 -346
rect 41146 -582 41382 -346
rect 40826 -902 41062 -666
rect 41146 -902 41382 -666
rect 38266 -5382 38502 -5146
rect 38586 -5382 38822 -5146
rect 38266 -5702 38502 -5466
rect 38586 -5702 38822 -5466
rect 31986 -6342 32222 -6106
rect 32306 -6342 32542 -6106
rect 31986 -6662 32222 -6426
rect 32306 -6662 32542 -6426
rect 44546 6938 44782 7174
rect 44866 6938 45102 7174
rect 44546 6618 44782 6854
rect 44866 6618 45102 6854
rect 44546 -2502 44782 -2266
rect 44866 -2502 45102 -2266
rect 44546 -2822 44782 -2586
rect 44866 -2822 45102 -2586
rect 48266 10658 48502 10894
rect 48586 10658 48822 10894
rect 48266 10338 48502 10574
rect 48586 10338 48822 10574
rect 50826 -1542 51062 -1306
rect 51146 -1542 51382 -1306
rect 50826 -1862 51062 -1626
rect 51146 -1862 51382 -1626
rect 51986 14378 52222 14614
rect 52306 14378 52542 14614
rect 51986 14058 52222 14294
rect 52306 14058 52542 14294
rect 48266 -4422 48502 -4186
rect 48586 -4422 48822 -4186
rect 48266 -4742 48502 -4506
rect 48586 -4742 48822 -4506
rect 41986 -7302 42222 -7066
rect 42306 -7302 42542 -7066
rect 41986 -7622 42222 -7386
rect 42306 -7622 42542 -7386
rect 54546 -3462 54782 -3226
rect 54866 -3462 55102 -3226
rect 54546 -3782 54782 -3546
rect 54866 -3782 55102 -3546
rect 60826 3218 61062 3454
rect 61146 3218 61382 3454
rect 60826 2898 61062 3134
rect 61146 2898 61382 3134
rect 60826 -582 61062 -346
rect 61146 -582 61382 -346
rect 60826 -902 61062 -666
rect 61146 -902 61382 -666
rect 58266 -5382 58502 -5146
rect 58586 -5382 58822 -5146
rect 58266 -5702 58502 -5466
rect 58586 -5702 58822 -5466
rect 51986 -6342 52222 -6106
rect 52306 -6342 52542 -6106
rect 51986 -6662 52222 -6426
rect 52306 -6662 52542 -6426
rect 64546 6938 64782 7174
rect 64866 6938 65102 7174
rect 64546 6618 64782 6854
rect 64866 6618 65102 6854
rect 64546 -2502 64782 -2266
rect 64866 -2502 65102 -2266
rect 64546 -2822 64782 -2586
rect 64866 -2822 65102 -2586
rect 68266 10658 68502 10894
rect 68586 10658 68822 10894
rect 68266 10338 68502 10574
rect 68586 10338 68822 10574
rect 70826 -1542 71062 -1306
rect 71146 -1542 71382 -1306
rect 70826 -1862 71062 -1626
rect 71146 -1862 71382 -1626
rect 71986 14378 72222 14614
rect 72306 14378 72542 14614
rect 71986 14058 72222 14294
rect 72306 14058 72542 14294
rect 68266 -4422 68502 -4186
rect 68586 -4422 68822 -4186
rect 68266 -4742 68502 -4506
rect 68586 -4742 68822 -4506
rect 61986 -7302 62222 -7066
rect 62306 -7302 62542 -7066
rect 61986 -7622 62222 -7386
rect 62306 -7622 62542 -7386
rect 74546 -3462 74782 -3226
rect 74866 -3462 75102 -3226
rect 74546 -3782 74782 -3546
rect 74866 -3782 75102 -3546
rect 78266 676658 78502 676894
rect 78586 676658 78822 676894
rect 78266 676338 78502 676574
rect 78586 676338 78822 676574
rect 78266 640658 78502 640894
rect 78586 640658 78822 640894
rect 78266 640338 78502 640574
rect 78586 640338 78822 640574
rect 78266 604658 78502 604894
rect 78586 604658 78822 604894
rect 78266 604338 78502 604574
rect 78586 604338 78822 604574
rect 78266 568658 78502 568894
rect 78586 568658 78822 568894
rect 78266 568338 78502 568574
rect 78586 568338 78822 568574
rect 78266 532658 78502 532894
rect 78586 532658 78822 532894
rect 78266 532338 78502 532574
rect 78586 532338 78822 532574
rect 78266 496658 78502 496894
rect 78586 496658 78822 496894
rect 78266 496338 78502 496574
rect 78586 496338 78822 496574
rect 78266 460658 78502 460894
rect 78586 460658 78822 460894
rect 78266 460338 78502 460574
rect 78586 460338 78822 460574
rect 78266 424658 78502 424894
rect 78586 424658 78822 424894
rect 78266 424338 78502 424574
rect 78586 424338 78822 424574
rect 78266 388658 78502 388894
rect 78586 388658 78822 388894
rect 78266 388338 78502 388574
rect 78586 388338 78822 388574
rect 78266 352658 78502 352894
rect 78586 352658 78822 352894
rect 78266 352338 78502 352574
rect 78586 352338 78822 352574
rect 78266 316658 78502 316894
rect 78586 316658 78822 316894
rect 78266 316338 78502 316574
rect 78586 316338 78822 316574
rect 78266 280658 78502 280894
rect 78586 280658 78822 280894
rect 78266 280338 78502 280574
rect 78586 280338 78822 280574
rect 78266 244658 78502 244894
rect 78586 244658 78822 244894
rect 78266 244338 78502 244574
rect 78586 244338 78822 244574
rect 78266 208658 78502 208894
rect 78586 208658 78822 208894
rect 78266 208338 78502 208574
rect 78586 208338 78822 208574
rect 78266 172658 78502 172894
rect 78586 172658 78822 172894
rect 78266 172338 78502 172574
rect 78586 172338 78822 172574
rect 78266 136658 78502 136894
rect 78586 136658 78822 136894
rect 78266 136338 78502 136574
rect 78586 136338 78822 136574
rect 78266 100658 78502 100894
rect 78586 100658 78822 100894
rect 78266 100338 78502 100574
rect 78586 100338 78822 100574
rect 78266 64658 78502 64894
rect 78586 64658 78822 64894
rect 78266 64338 78502 64574
rect 78586 64338 78822 64574
rect 78266 28658 78502 28894
rect 78586 28658 78822 28894
rect 78266 28338 78502 28574
rect 78586 28338 78822 28574
rect 80826 704602 81062 704838
rect 81146 704602 81382 704838
rect 80826 704282 81062 704518
rect 81146 704282 81382 704518
rect 80826 687218 81062 687454
rect 81146 687218 81382 687454
rect 80826 686898 81062 687134
rect 81146 686898 81382 687134
rect 80826 651218 81062 651454
rect 81146 651218 81382 651454
rect 80826 650898 81062 651134
rect 81146 650898 81382 651134
rect 80826 615218 81062 615454
rect 81146 615218 81382 615454
rect 80826 614898 81062 615134
rect 81146 614898 81382 615134
rect 80826 579218 81062 579454
rect 81146 579218 81382 579454
rect 80826 578898 81062 579134
rect 81146 578898 81382 579134
rect 80826 543218 81062 543454
rect 81146 543218 81382 543454
rect 80826 542898 81062 543134
rect 81146 542898 81382 543134
rect 80826 507218 81062 507454
rect 81146 507218 81382 507454
rect 80826 506898 81062 507134
rect 81146 506898 81382 507134
rect 80826 471218 81062 471454
rect 81146 471218 81382 471454
rect 80826 470898 81062 471134
rect 81146 470898 81382 471134
rect 80826 435218 81062 435454
rect 81146 435218 81382 435454
rect 80826 434898 81062 435134
rect 81146 434898 81382 435134
rect 80826 399218 81062 399454
rect 81146 399218 81382 399454
rect 80826 398898 81062 399134
rect 81146 398898 81382 399134
rect 80826 363218 81062 363454
rect 81146 363218 81382 363454
rect 80826 362898 81062 363134
rect 81146 362898 81382 363134
rect 80826 327218 81062 327454
rect 81146 327218 81382 327454
rect 80826 326898 81062 327134
rect 81146 326898 81382 327134
rect 80826 291218 81062 291454
rect 81146 291218 81382 291454
rect 80826 290898 81062 291134
rect 81146 290898 81382 291134
rect 80826 255218 81062 255454
rect 81146 255218 81382 255454
rect 80826 254898 81062 255134
rect 81146 254898 81382 255134
rect 80826 219218 81062 219454
rect 81146 219218 81382 219454
rect 80826 218898 81062 219134
rect 81146 218898 81382 219134
rect 80826 183218 81062 183454
rect 81146 183218 81382 183454
rect 80826 182898 81062 183134
rect 81146 182898 81382 183134
rect 80826 147218 81062 147454
rect 81146 147218 81382 147454
rect 80826 146898 81062 147134
rect 81146 146898 81382 147134
rect 80826 111218 81062 111454
rect 81146 111218 81382 111454
rect 80826 110898 81062 111134
rect 81146 110898 81382 111134
rect 80826 75218 81062 75454
rect 81146 75218 81382 75454
rect 80826 74898 81062 75134
rect 81146 74898 81382 75134
rect 80826 39218 81062 39454
rect 81146 39218 81382 39454
rect 80826 38898 81062 39134
rect 81146 38898 81382 39134
rect 80826 3218 81062 3454
rect 81146 3218 81382 3454
rect 80826 2898 81062 3134
rect 81146 2898 81382 3134
rect 80826 -582 81062 -346
rect 81146 -582 81382 -346
rect 80826 -902 81062 -666
rect 81146 -902 81382 -666
rect 91986 710362 92222 710598
rect 92306 710362 92542 710598
rect 91986 710042 92222 710278
rect 92306 710042 92542 710278
rect 88266 708442 88502 708678
rect 88586 708442 88822 708678
rect 88266 708122 88502 708358
rect 88586 708122 88822 708358
rect 81986 680378 82222 680614
rect 82306 680378 82542 680614
rect 81986 680058 82222 680294
rect 82306 680058 82542 680294
rect 81986 644378 82222 644614
rect 82306 644378 82542 644614
rect 81986 644058 82222 644294
rect 82306 644058 82542 644294
rect 81986 608378 82222 608614
rect 82306 608378 82542 608614
rect 81986 608058 82222 608294
rect 82306 608058 82542 608294
rect 81986 572378 82222 572614
rect 82306 572378 82542 572614
rect 81986 572058 82222 572294
rect 82306 572058 82542 572294
rect 81986 536378 82222 536614
rect 82306 536378 82542 536614
rect 81986 536058 82222 536294
rect 82306 536058 82542 536294
rect 81986 500378 82222 500614
rect 82306 500378 82542 500614
rect 81986 500058 82222 500294
rect 82306 500058 82542 500294
rect 81986 464378 82222 464614
rect 82306 464378 82542 464614
rect 81986 464058 82222 464294
rect 82306 464058 82542 464294
rect 81986 428378 82222 428614
rect 82306 428378 82542 428614
rect 81986 428058 82222 428294
rect 82306 428058 82542 428294
rect 81986 392378 82222 392614
rect 82306 392378 82542 392614
rect 81986 392058 82222 392294
rect 82306 392058 82542 392294
rect 81986 356378 82222 356614
rect 82306 356378 82542 356614
rect 81986 356058 82222 356294
rect 82306 356058 82542 356294
rect 81986 320378 82222 320614
rect 82306 320378 82542 320614
rect 81986 320058 82222 320294
rect 82306 320058 82542 320294
rect 81986 284378 82222 284614
rect 82306 284378 82542 284614
rect 81986 284058 82222 284294
rect 82306 284058 82542 284294
rect 81986 248378 82222 248614
rect 82306 248378 82542 248614
rect 81986 248058 82222 248294
rect 82306 248058 82542 248294
rect 81986 212378 82222 212614
rect 82306 212378 82542 212614
rect 81986 212058 82222 212294
rect 82306 212058 82542 212294
rect 81986 176378 82222 176614
rect 82306 176378 82542 176614
rect 81986 176058 82222 176294
rect 82306 176058 82542 176294
rect 81986 140378 82222 140614
rect 82306 140378 82542 140614
rect 81986 140058 82222 140294
rect 82306 140058 82542 140294
rect 81986 104378 82222 104614
rect 82306 104378 82542 104614
rect 81986 104058 82222 104294
rect 82306 104058 82542 104294
rect 81986 68378 82222 68614
rect 82306 68378 82542 68614
rect 81986 68058 82222 68294
rect 82306 68058 82542 68294
rect 81986 32378 82222 32614
rect 82306 32378 82542 32614
rect 81986 32058 82222 32294
rect 82306 32058 82542 32294
rect 78266 -5382 78502 -5146
rect 78586 -5382 78822 -5146
rect 78266 -5702 78502 -5466
rect 78586 -5702 78822 -5466
rect 71986 -6342 72222 -6106
rect 72306 -6342 72542 -6106
rect 71986 -6662 72222 -6426
rect 72306 -6662 72542 -6426
rect 84546 706522 84782 706758
rect 84866 706522 85102 706758
rect 84546 706202 84782 706438
rect 84866 706202 85102 706438
rect 84546 690938 84782 691174
rect 84866 690938 85102 691174
rect 84546 690618 84782 690854
rect 84866 690618 85102 690854
rect 84546 654938 84782 655174
rect 84866 654938 85102 655174
rect 84546 654618 84782 654854
rect 84866 654618 85102 654854
rect 84546 618938 84782 619174
rect 84866 618938 85102 619174
rect 84546 618618 84782 618854
rect 84866 618618 85102 618854
rect 84546 582938 84782 583174
rect 84866 582938 85102 583174
rect 84546 582618 84782 582854
rect 84866 582618 85102 582854
rect 84546 546938 84782 547174
rect 84866 546938 85102 547174
rect 84546 546618 84782 546854
rect 84866 546618 85102 546854
rect 84546 510938 84782 511174
rect 84866 510938 85102 511174
rect 84546 510618 84782 510854
rect 84866 510618 85102 510854
rect 84546 474938 84782 475174
rect 84866 474938 85102 475174
rect 84546 474618 84782 474854
rect 84866 474618 85102 474854
rect 84546 438938 84782 439174
rect 84866 438938 85102 439174
rect 84546 438618 84782 438854
rect 84866 438618 85102 438854
rect 84546 402938 84782 403174
rect 84866 402938 85102 403174
rect 84546 402618 84782 402854
rect 84866 402618 85102 402854
rect 84546 366938 84782 367174
rect 84866 366938 85102 367174
rect 84546 366618 84782 366854
rect 84866 366618 85102 366854
rect 84546 330938 84782 331174
rect 84866 330938 85102 331174
rect 84546 330618 84782 330854
rect 84866 330618 85102 330854
rect 84546 294938 84782 295174
rect 84866 294938 85102 295174
rect 84546 294618 84782 294854
rect 84866 294618 85102 294854
rect 84546 258938 84782 259174
rect 84866 258938 85102 259174
rect 84546 258618 84782 258854
rect 84866 258618 85102 258854
rect 84546 222938 84782 223174
rect 84866 222938 85102 223174
rect 84546 222618 84782 222854
rect 84866 222618 85102 222854
rect 84546 186938 84782 187174
rect 84866 186938 85102 187174
rect 84546 186618 84782 186854
rect 84866 186618 85102 186854
rect 84546 150938 84782 151174
rect 84866 150938 85102 151174
rect 84546 150618 84782 150854
rect 84866 150618 85102 150854
rect 84546 114938 84782 115174
rect 84866 114938 85102 115174
rect 84546 114618 84782 114854
rect 84866 114618 85102 114854
rect 84546 78938 84782 79174
rect 84866 78938 85102 79174
rect 84546 78618 84782 78854
rect 84866 78618 85102 78854
rect 84546 42938 84782 43174
rect 84866 42938 85102 43174
rect 84546 42618 84782 42854
rect 84866 42618 85102 42854
rect 84546 6938 84782 7174
rect 84866 6938 85102 7174
rect 84546 6618 84782 6854
rect 84866 6618 85102 6854
rect 84546 -2502 84782 -2266
rect 84866 -2502 85102 -2266
rect 84546 -2822 84782 -2586
rect 84866 -2822 85102 -2586
rect 88266 694658 88502 694894
rect 88586 694658 88822 694894
rect 88266 694338 88502 694574
rect 88586 694338 88822 694574
rect 88266 658658 88502 658894
rect 88586 658658 88822 658894
rect 88266 658338 88502 658574
rect 88586 658338 88822 658574
rect 88266 622658 88502 622894
rect 88586 622658 88822 622894
rect 88266 622338 88502 622574
rect 88586 622338 88822 622574
rect 88266 586658 88502 586894
rect 88586 586658 88822 586894
rect 88266 586338 88502 586574
rect 88586 586338 88822 586574
rect 88266 550658 88502 550894
rect 88586 550658 88822 550894
rect 88266 550338 88502 550574
rect 88586 550338 88822 550574
rect 88266 514658 88502 514894
rect 88586 514658 88822 514894
rect 88266 514338 88502 514574
rect 88586 514338 88822 514574
rect 88266 478658 88502 478894
rect 88586 478658 88822 478894
rect 88266 478338 88502 478574
rect 88586 478338 88822 478574
rect 88266 442658 88502 442894
rect 88586 442658 88822 442894
rect 88266 442338 88502 442574
rect 88586 442338 88822 442574
rect 88266 406658 88502 406894
rect 88586 406658 88822 406894
rect 88266 406338 88502 406574
rect 88586 406338 88822 406574
rect 88266 370658 88502 370894
rect 88586 370658 88822 370894
rect 88266 370338 88502 370574
rect 88586 370338 88822 370574
rect 88266 334658 88502 334894
rect 88586 334658 88822 334894
rect 88266 334338 88502 334574
rect 88586 334338 88822 334574
rect 88266 298658 88502 298894
rect 88586 298658 88822 298894
rect 88266 298338 88502 298574
rect 88586 298338 88822 298574
rect 88266 262658 88502 262894
rect 88586 262658 88822 262894
rect 88266 262338 88502 262574
rect 88586 262338 88822 262574
rect 88266 226658 88502 226894
rect 88586 226658 88822 226894
rect 88266 226338 88502 226574
rect 88586 226338 88822 226574
rect 88266 190658 88502 190894
rect 88586 190658 88822 190894
rect 88266 190338 88502 190574
rect 88586 190338 88822 190574
rect 88266 154658 88502 154894
rect 88586 154658 88822 154894
rect 88266 154338 88502 154574
rect 88586 154338 88822 154574
rect 88266 118658 88502 118894
rect 88586 118658 88822 118894
rect 88266 118338 88502 118574
rect 88586 118338 88822 118574
rect 88266 82658 88502 82894
rect 88586 82658 88822 82894
rect 88266 82338 88502 82574
rect 88586 82338 88822 82574
rect 88266 46658 88502 46894
rect 88586 46658 88822 46894
rect 88266 46338 88502 46574
rect 88586 46338 88822 46574
rect 88266 10658 88502 10894
rect 88586 10658 88822 10894
rect 88266 10338 88502 10574
rect 88586 10338 88822 10574
rect 90826 705562 91062 705798
rect 91146 705562 91382 705798
rect 90826 705242 91062 705478
rect 91146 705242 91382 705478
rect 90826 669218 91062 669454
rect 91146 669218 91382 669454
rect 90826 668898 91062 669134
rect 91146 668898 91382 669134
rect 90826 633218 91062 633454
rect 91146 633218 91382 633454
rect 90826 632898 91062 633134
rect 91146 632898 91382 633134
rect 90826 597218 91062 597454
rect 91146 597218 91382 597454
rect 90826 596898 91062 597134
rect 91146 596898 91382 597134
rect 90826 561218 91062 561454
rect 91146 561218 91382 561454
rect 90826 560898 91062 561134
rect 91146 560898 91382 561134
rect 90826 525218 91062 525454
rect 91146 525218 91382 525454
rect 90826 524898 91062 525134
rect 91146 524898 91382 525134
rect 90826 489218 91062 489454
rect 91146 489218 91382 489454
rect 90826 488898 91062 489134
rect 91146 488898 91382 489134
rect 90826 453218 91062 453454
rect 91146 453218 91382 453454
rect 90826 452898 91062 453134
rect 91146 452898 91382 453134
rect 90826 417218 91062 417454
rect 91146 417218 91382 417454
rect 90826 416898 91062 417134
rect 91146 416898 91382 417134
rect 90826 381218 91062 381454
rect 91146 381218 91382 381454
rect 90826 380898 91062 381134
rect 91146 380898 91382 381134
rect 90826 345218 91062 345454
rect 91146 345218 91382 345454
rect 90826 344898 91062 345134
rect 91146 344898 91382 345134
rect 90826 309218 91062 309454
rect 91146 309218 91382 309454
rect 90826 308898 91062 309134
rect 91146 308898 91382 309134
rect 90826 273218 91062 273454
rect 91146 273218 91382 273454
rect 90826 272898 91062 273134
rect 91146 272898 91382 273134
rect 90826 237218 91062 237454
rect 91146 237218 91382 237454
rect 90826 236898 91062 237134
rect 91146 236898 91382 237134
rect 90826 201218 91062 201454
rect 91146 201218 91382 201454
rect 90826 200898 91062 201134
rect 91146 200898 91382 201134
rect 90826 165218 91062 165454
rect 91146 165218 91382 165454
rect 90826 164898 91062 165134
rect 91146 164898 91382 165134
rect 90826 129218 91062 129454
rect 91146 129218 91382 129454
rect 90826 128898 91062 129134
rect 91146 128898 91382 129134
rect 90826 93218 91062 93454
rect 91146 93218 91382 93454
rect 90826 92898 91062 93134
rect 91146 92898 91382 93134
rect 90826 57218 91062 57454
rect 91146 57218 91382 57454
rect 90826 56898 91062 57134
rect 91146 56898 91382 57134
rect 90826 21218 91062 21454
rect 91146 21218 91382 21454
rect 90826 20898 91062 21134
rect 91146 20898 91382 21134
rect 90826 -1542 91062 -1306
rect 91146 -1542 91382 -1306
rect 90826 -1862 91062 -1626
rect 91146 -1862 91382 -1626
rect 101986 711322 102222 711558
rect 102306 711322 102542 711558
rect 101986 711002 102222 711238
rect 102306 711002 102542 711238
rect 98266 709402 98502 709638
rect 98586 709402 98822 709638
rect 98266 709082 98502 709318
rect 98586 709082 98822 709318
rect 91986 698378 92222 698614
rect 92306 698378 92542 698614
rect 91986 698058 92222 698294
rect 92306 698058 92542 698294
rect 91986 662378 92222 662614
rect 92306 662378 92542 662614
rect 91986 662058 92222 662294
rect 92306 662058 92542 662294
rect 91986 626378 92222 626614
rect 92306 626378 92542 626614
rect 91986 626058 92222 626294
rect 92306 626058 92542 626294
rect 91986 590378 92222 590614
rect 92306 590378 92542 590614
rect 91986 590058 92222 590294
rect 92306 590058 92542 590294
rect 91986 554378 92222 554614
rect 92306 554378 92542 554614
rect 91986 554058 92222 554294
rect 92306 554058 92542 554294
rect 91986 518378 92222 518614
rect 92306 518378 92542 518614
rect 91986 518058 92222 518294
rect 92306 518058 92542 518294
rect 91986 482378 92222 482614
rect 92306 482378 92542 482614
rect 91986 482058 92222 482294
rect 92306 482058 92542 482294
rect 91986 446378 92222 446614
rect 92306 446378 92542 446614
rect 91986 446058 92222 446294
rect 92306 446058 92542 446294
rect 91986 410378 92222 410614
rect 92306 410378 92542 410614
rect 91986 410058 92222 410294
rect 92306 410058 92542 410294
rect 91986 374378 92222 374614
rect 92306 374378 92542 374614
rect 91986 374058 92222 374294
rect 92306 374058 92542 374294
rect 91986 338378 92222 338614
rect 92306 338378 92542 338614
rect 91986 338058 92222 338294
rect 92306 338058 92542 338294
rect 91986 302378 92222 302614
rect 92306 302378 92542 302614
rect 91986 302058 92222 302294
rect 92306 302058 92542 302294
rect 91986 266378 92222 266614
rect 92306 266378 92542 266614
rect 91986 266058 92222 266294
rect 92306 266058 92542 266294
rect 91986 230378 92222 230614
rect 92306 230378 92542 230614
rect 91986 230058 92222 230294
rect 92306 230058 92542 230294
rect 91986 194378 92222 194614
rect 92306 194378 92542 194614
rect 91986 194058 92222 194294
rect 92306 194058 92542 194294
rect 91986 158378 92222 158614
rect 92306 158378 92542 158614
rect 91986 158058 92222 158294
rect 92306 158058 92542 158294
rect 91986 122378 92222 122614
rect 92306 122378 92542 122614
rect 91986 122058 92222 122294
rect 92306 122058 92542 122294
rect 91986 86378 92222 86614
rect 92306 86378 92542 86614
rect 91986 86058 92222 86294
rect 92306 86058 92542 86294
rect 91986 50378 92222 50614
rect 92306 50378 92542 50614
rect 91986 50058 92222 50294
rect 92306 50058 92542 50294
rect 91986 14378 92222 14614
rect 92306 14378 92542 14614
rect 91986 14058 92222 14294
rect 92306 14058 92542 14294
rect 88266 -4422 88502 -4186
rect 88586 -4422 88822 -4186
rect 88266 -4742 88502 -4506
rect 88586 -4742 88822 -4506
rect 81986 -7302 82222 -7066
rect 82306 -7302 82542 -7066
rect 81986 -7622 82222 -7386
rect 82306 -7622 82542 -7386
rect 94546 707482 94782 707718
rect 94866 707482 95102 707718
rect 94546 707162 94782 707398
rect 94866 707162 95102 707398
rect 94546 672938 94782 673174
rect 94866 672938 95102 673174
rect 94546 672618 94782 672854
rect 94866 672618 95102 672854
rect 94546 636938 94782 637174
rect 94866 636938 95102 637174
rect 94546 636618 94782 636854
rect 94866 636618 95102 636854
rect 94546 600938 94782 601174
rect 94866 600938 95102 601174
rect 94546 600618 94782 600854
rect 94866 600618 95102 600854
rect 94546 564938 94782 565174
rect 94866 564938 95102 565174
rect 94546 564618 94782 564854
rect 94866 564618 95102 564854
rect 94546 528938 94782 529174
rect 94866 528938 95102 529174
rect 94546 528618 94782 528854
rect 94866 528618 95102 528854
rect 94546 492938 94782 493174
rect 94866 492938 95102 493174
rect 94546 492618 94782 492854
rect 94866 492618 95102 492854
rect 94546 456938 94782 457174
rect 94866 456938 95102 457174
rect 94546 456618 94782 456854
rect 94866 456618 95102 456854
rect 94546 420938 94782 421174
rect 94866 420938 95102 421174
rect 94546 420618 94782 420854
rect 94866 420618 95102 420854
rect 94546 384938 94782 385174
rect 94866 384938 95102 385174
rect 94546 384618 94782 384854
rect 94866 384618 95102 384854
rect 94546 348938 94782 349174
rect 94866 348938 95102 349174
rect 94546 348618 94782 348854
rect 94866 348618 95102 348854
rect 94546 312938 94782 313174
rect 94866 312938 95102 313174
rect 94546 312618 94782 312854
rect 94866 312618 95102 312854
rect 94546 276938 94782 277174
rect 94866 276938 95102 277174
rect 94546 276618 94782 276854
rect 94866 276618 95102 276854
rect 94546 240938 94782 241174
rect 94866 240938 95102 241174
rect 94546 240618 94782 240854
rect 94866 240618 95102 240854
rect 94546 204938 94782 205174
rect 94866 204938 95102 205174
rect 94546 204618 94782 204854
rect 94866 204618 95102 204854
rect 94546 168938 94782 169174
rect 94866 168938 95102 169174
rect 94546 168618 94782 168854
rect 94866 168618 95102 168854
rect 94546 132938 94782 133174
rect 94866 132938 95102 133174
rect 94546 132618 94782 132854
rect 94866 132618 95102 132854
rect 94546 96938 94782 97174
rect 94866 96938 95102 97174
rect 94546 96618 94782 96854
rect 94866 96618 95102 96854
rect 94546 60938 94782 61174
rect 94866 60938 95102 61174
rect 94546 60618 94782 60854
rect 94866 60618 95102 60854
rect 94546 24938 94782 25174
rect 94866 24938 95102 25174
rect 94546 24618 94782 24854
rect 94866 24618 95102 24854
rect 94546 -3462 94782 -3226
rect 94866 -3462 95102 -3226
rect 94546 -3782 94782 -3546
rect 94866 -3782 95102 -3546
rect 98266 676658 98502 676894
rect 98586 676658 98822 676894
rect 98266 676338 98502 676574
rect 98586 676338 98822 676574
rect 98266 640658 98502 640894
rect 98586 640658 98822 640894
rect 98266 640338 98502 640574
rect 98586 640338 98822 640574
rect 98266 604658 98502 604894
rect 98586 604658 98822 604894
rect 98266 604338 98502 604574
rect 98586 604338 98822 604574
rect 98266 568658 98502 568894
rect 98586 568658 98822 568894
rect 98266 568338 98502 568574
rect 98586 568338 98822 568574
rect 98266 532658 98502 532894
rect 98586 532658 98822 532894
rect 98266 532338 98502 532574
rect 98586 532338 98822 532574
rect 98266 496658 98502 496894
rect 98586 496658 98822 496894
rect 98266 496338 98502 496574
rect 98586 496338 98822 496574
rect 98266 460658 98502 460894
rect 98586 460658 98822 460894
rect 98266 460338 98502 460574
rect 98586 460338 98822 460574
rect 98266 424658 98502 424894
rect 98586 424658 98822 424894
rect 98266 424338 98502 424574
rect 98586 424338 98822 424574
rect 98266 388658 98502 388894
rect 98586 388658 98822 388894
rect 98266 388338 98502 388574
rect 98586 388338 98822 388574
rect 98266 352658 98502 352894
rect 98586 352658 98822 352894
rect 98266 352338 98502 352574
rect 98586 352338 98822 352574
rect 98266 316658 98502 316894
rect 98586 316658 98822 316894
rect 98266 316338 98502 316574
rect 98586 316338 98822 316574
rect 98266 280658 98502 280894
rect 98586 280658 98822 280894
rect 98266 280338 98502 280574
rect 98586 280338 98822 280574
rect 98266 244658 98502 244894
rect 98586 244658 98822 244894
rect 98266 244338 98502 244574
rect 98586 244338 98822 244574
rect 98266 208658 98502 208894
rect 98586 208658 98822 208894
rect 98266 208338 98502 208574
rect 98586 208338 98822 208574
rect 98266 172658 98502 172894
rect 98586 172658 98822 172894
rect 98266 172338 98502 172574
rect 98586 172338 98822 172574
rect 98266 136658 98502 136894
rect 98586 136658 98822 136894
rect 98266 136338 98502 136574
rect 98586 136338 98822 136574
rect 98266 100658 98502 100894
rect 98586 100658 98822 100894
rect 98266 100338 98502 100574
rect 98586 100338 98822 100574
rect 98266 64658 98502 64894
rect 98586 64658 98822 64894
rect 98266 64338 98502 64574
rect 98586 64338 98822 64574
rect 98266 28658 98502 28894
rect 98586 28658 98822 28894
rect 98266 28338 98502 28574
rect 98586 28338 98822 28574
rect 100826 704602 101062 704838
rect 101146 704602 101382 704838
rect 100826 704282 101062 704518
rect 101146 704282 101382 704518
rect 100826 687218 101062 687454
rect 101146 687218 101382 687454
rect 100826 686898 101062 687134
rect 101146 686898 101382 687134
rect 100826 651218 101062 651454
rect 101146 651218 101382 651454
rect 100826 650898 101062 651134
rect 101146 650898 101382 651134
rect 100826 615218 101062 615454
rect 101146 615218 101382 615454
rect 100826 614898 101062 615134
rect 101146 614898 101382 615134
rect 100826 579218 101062 579454
rect 101146 579218 101382 579454
rect 100826 578898 101062 579134
rect 101146 578898 101382 579134
rect 100826 543218 101062 543454
rect 101146 543218 101382 543454
rect 100826 542898 101062 543134
rect 101146 542898 101382 543134
rect 100826 507218 101062 507454
rect 101146 507218 101382 507454
rect 100826 506898 101062 507134
rect 101146 506898 101382 507134
rect 100826 471218 101062 471454
rect 101146 471218 101382 471454
rect 100826 470898 101062 471134
rect 101146 470898 101382 471134
rect 100826 435218 101062 435454
rect 101146 435218 101382 435454
rect 100826 434898 101062 435134
rect 101146 434898 101382 435134
rect 100826 399218 101062 399454
rect 101146 399218 101382 399454
rect 100826 398898 101062 399134
rect 101146 398898 101382 399134
rect 100826 363218 101062 363454
rect 101146 363218 101382 363454
rect 100826 362898 101062 363134
rect 101146 362898 101382 363134
rect 100826 327218 101062 327454
rect 101146 327218 101382 327454
rect 100826 326898 101062 327134
rect 101146 326898 101382 327134
rect 100826 291218 101062 291454
rect 101146 291218 101382 291454
rect 100826 290898 101062 291134
rect 101146 290898 101382 291134
rect 100826 255218 101062 255454
rect 101146 255218 101382 255454
rect 100826 254898 101062 255134
rect 101146 254898 101382 255134
rect 100826 219218 101062 219454
rect 101146 219218 101382 219454
rect 100826 218898 101062 219134
rect 101146 218898 101382 219134
rect 100826 183218 101062 183454
rect 101146 183218 101382 183454
rect 100826 182898 101062 183134
rect 101146 182898 101382 183134
rect 100826 147218 101062 147454
rect 101146 147218 101382 147454
rect 100826 146898 101062 147134
rect 101146 146898 101382 147134
rect 100826 111218 101062 111454
rect 101146 111218 101382 111454
rect 100826 110898 101062 111134
rect 101146 110898 101382 111134
rect 100826 75218 101062 75454
rect 101146 75218 101382 75454
rect 100826 74898 101062 75134
rect 101146 74898 101382 75134
rect 100826 39218 101062 39454
rect 101146 39218 101382 39454
rect 100826 38898 101062 39134
rect 101146 38898 101382 39134
rect 100826 3218 101062 3454
rect 101146 3218 101382 3454
rect 100826 2898 101062 3134
rect 101146 2898 101382 3134
rect 100826 -582 101062 -346
rect 101146 -582 101382 -346
rect 100826 -902 101062 -666
rect 101146 -902 101382 -666
rect 111986 710362 112222 710598
rect 112306 710362 112542 710598
rect 111986 710042 112222 710278
rect 112306 710042 112542 710278
rect 108266 708442 108502 708678
rect 108586 708442 108822 708678
rect 108266 708122 108502 708358
rect 108586 708122 108822 708358
rect 101986 680378 102222 680614
rect 102306 680378 102542 680614
rect 101986 680058 102222 680294
rect 102306 680058 102542 680294
rect 101986 644378 102222 644614
rect 102306 644378 102542 644614
rect 101986 644058 102222 644294
rect 102306 644058 102542 644294
rect 101986 608378 102222 608614
rect 102306 608378 102542 608614
rect 101986 608058 102222 608294
rect 102306 608058 102542 608294
rect 101986 572378 102222 572614
rect 102306 572378 102542 572614
rect 101986 572058 102222 572294
rect 102306 572058 102542 572294
rect 101986 536378 102222 536614
rect 102306 536378 102542 536614
rect 101986 536058 102222 536294
rect 102306 536058 102542 536294
rect 101986 500378 102222 500614
rect 102306 500378 102542 500614
rect 101986 500058 102222 500294
rect 102306 500058 102542 500294
rect 101986 464378 102222 464614
rect 102306 464378 102542 464614
rect 101986 464058 102222 464294
rect 102306 464058 102542 464294
rect 101986 428378 102222 428614
rect 102306 428378 102542 428614
rect 101986 428058 102222 428294
rect 102306 428058 102542 428294
rect 101986 392378 102222 392614
rect 102306 392378 102542 392614
rect 101986 392058 102222 392294
rect 102306 392058 102542 392294
rect 101986 356378 102222 356614
rect 102306 356378 102542 356614
rect 101986 356058 102222 356294
rect 102306 356058 102542 356294
rect 101986 320378 102222 320614
rect 102306 320378 102542 320614
rect 101986 320058 102222 320294
rect 102306 320058 102542 320294
rect 101986 284378 102222 284614
rect 102306 284378 102542 284614
rect 101986 284058 102222 284294
rect 102306 284058 102542 284294
rect 101986 248378 102222 248614
rect 102306 248378 102542 248614
rect 101986 248058 102222 248294
rect 102306 248058 102542 248294
rect 101986 212378 102222 212614
rect 102306 212378 102542 212614
rect 101986 212058 102222 212294
rect 102306 212058 102542 212294
rect 101986 176378 102222 176614
rect 102306 176378 102542 176614
rect 101986 176058 102222 176294
rect 102306 176058 102542 176294
rect 101986 140378 102222 140614
rect 102306 140378 102542 140614
rect 101986 140058 102222 140294
rect 102306 140058 102542 140294
rect 101986 104378 102222 104614
rect 102306 104378 102542 104614
rect 101986 104058 102222 104294
rect 102306 104058 102542 104294
rect 101986 68378 102222 68614
rect 102306 68378 102542 68614
rect 101986 68058 102222 68294
rect 102306 68058 102542 68294
rect 101986 32378 102222 32614
rect 102306 32378 102542 32614
rect 101986 32058 102222 32294
rect 102306 32058 102542 32294
rect 98266 -5382 98502 -5146
rect 98586 -5382 98822 -5146
rect 98266 -5702 98502 -5466
rect 98586 -5702 98822 -5466
rect 91986 -6342 92222 -6106
rect 92306 -6342 92542 -6106
rect 91986 -6662 92222 -6426
rect 92306 -6662 92542 -6426
rect 104546 706522 104782 706758
rect 104866 706522 105102 706758
rect 104546 706202 104782 706438
rect 104866 706202 105102 706438
rect 104546 690938 104782 691174
rect 104866 690938 105102 691174
rect 104546 690618 104782 690854
rect 104866 690618 105102 690854
rect 104546 654938 104782 655174
rect 104866 654938 105102 655174
rect 104546 654618 104782 654854
rect 104866 654618 105102 654854
rect 104546 618938 104782 619174
rect 104866 618938 105102 619174
rect 104546 618618 104782 618854
rect 104866 618618 105102 618854
rect 104546 582938 104782 583174
rect 104866 582938 105102 583174
rect 104546 582618 104782 582854
rect 104866 582618 105102 582854
rect 104546 546938 104782 547174
rect 104866 546938 105102 547174
rect 104546 546618 104782 546854
rect 104866 546618 105102 546854
rect 104546 510938 104782 511174
rect 104866 510938 105102 511174
rect 104546 510618 104782 510854
rect 104866 510618 105102 510854
rect 104546 474938 104782 475174
rect 104866 474938 105102 475174
rect 104546 474618 104782 474854
rect 104866 474618 105102 474854
rect 104546 438938 104782 439174
rect 104866 438938 105102 439174
rect 104546 438618 104782 438854
rect 104866 438618 105102 438854
rect 104546 402938 104782 403174
rect 104866 402938 105102 403174
rect 104546 402618 104782 402854
rect 104866 402618 105102 402854
rect 104546 366938 104782 367174
rect 104866 366938 105102 367174
rect 104546 366618 104782 366854
rect 104866 366618 105102 366854
rect 104546 330938 104782 331174
rect 104866 330938 105102 331174
rect 104546 330618 104782 330854
rect 104866 330618 105102 330854
rect 104546 294938 104782 295174
rect 104866 294938 105102 295174
rect 104546 294618 104782 294854
rect 104866 294618 105102 294854
rect 104546 258938 104782 259174
rect 104866 258938 105102 259174
rect 104546 258618 104782 258854
rect 104866 258618 105102 258854
rect 104546 222938 104782 223174
rect 104866 222938 105102 223174
rect 104546 222618 104782 222854
rect 104866 222618 105102 222854
rect 104546 186938 104782 187174
rect 104866 186938 105102 187174
rect 104546 186618 104782 186854
rect 104866 186618 105102 186854
rect 104546 150938 104782 151174
rect 104866 150938 105102 151174
rect 104546 150618 104782 150854
rect 104866 150618 105102 150854
rect 104546 114938 104782 115174
rect 104866 114938 105102 115174
rect 104546 114618 104782 114854
rect 104866 114618 105102 114854
rect 104546 78938 104782 79174
rect 104866 78938 105102 79174
rect 104546 78618 104782 78854
rect 104866 78618 105102 78854
rect 104546 42938 104782 43174
rect 104866 42938 105102 43174
rect 104546 42618 104782 42854
rect 104866 42618 105102 42854
rect 104546 6938 104782 7174
rect 104866 6938 105102 7174
rect 104546 6618 104782 6854
rect 104866 6618 105102 6854
rect 104546 -2502 104782 -2266
rect 104866 -2502 105102 -2266
rect 104546 -2822 104782 -2586
rect 104866 -2822 105102 -2586
rect 108266 694658 108502 694894
rect 108586 694658 108822 694894
rect 108266 694338 108502 694574
rect 108586 694338 108822 694574
rect 108266 658658 108502 658894
rect 108586 658658 108822 658894
rect 108266 658338 108502 658574
rect 108586 658338 108822 658574
rect 108266 622658 108502 622894
rect 108586 622658 108822 622894
rect 108266 622338 108502 622574
rect 108586 622338 108822 622574
rect 108266 586658 108502 586894
rect 108586 586658 108822 586894
rect 108266 586338 108502 586574
rect 108586 586338 108822 586574
rect 108266 550658 108502 550894
rect 108586 550658 108822 550894
rect 108266 550338 108502 550574
rect 108586 550338 108822 550574
rect 108266 514658 108502 514894
rect 108586 514658 108822 514894
rect 108266 514338 108502 514574
rect 108586 514338 108822 514574
rect 108266 478658 108502 478894
rect 108586 478658 108822 478894
rect 108266 478338 108502 478574
rect 108586 478338 108822 478574
rect 108266 442658 108502 442894
rect 108586 442658 108822 442894
rect 108266 442338 108502 442574
rect 108586 442338 108822 442574
rect 108266 406658 108502 406894
rect 108586 406658 108822 406894
rect 108266 406338 108502 406574
rect 108586 406338 108822 406574
rect 108266 370658 108502 370894
rect 108586 370658 108822 370894
rect 108266 370338 108502 370574
rect 108586 370338 108822 370574
rect 108266 334658 108502 334894
rect 108586 334658 108822 334894
rect 108266 334338 108502 334574
rect 108586 334338 108822 334574
rect 108266 298658 108502 298894
rect 108586 298658 108822 298894
rect 108266 298338 108502 298574
rect 108586 298338 108822 298574
rect 108266 262658 108502 262894
rect 108586 262658 108822 262894
rect 108266 262338 108502 262574
rect 108586 262338 108822 262574
rect 108266 226658 108502 226894
rect 108586 226658 108822 226894
rect 108266 226338 108502 226574
rect 108586 226338 108822 226574
rect 108266 190658 108502 190894
rect 108586 190658 108822 190894
rect 108266 190338 108502 190574
rect 108586 190338 108822 190574
rect 108266 154658 108502 154894
rect 108586 154658 108822 154894
rect 108266 154338 108502 154574
rect 108586 154338 108822 154574
rect 108266 118658 108502 118894
rect 108586 118658 108822 118894
rect 108266 118338 108502 118574
rect 108586 118338 108822 118574
rect 108266 82658 108502 82894
rect 108586 82658 108822 82894
rect 108266 82338 108502 82574
rect 108586 82338 108822 82574
rect 108266 46658 108502 46894
rect 108586 46658 108822 46894
rect 108266 46338 108502 46574
rect 108586 46338 108822 46574
rect 108266 10658 108502 10894
rect 108586 10658 108822 10894
rect 108266 10338 108502 10574
rect 108586 10338 108822 10574
rect 110826 705562 111062 705798
rect 111146 705562 111382 705798
rect 110826 705242 111062 705478
rect 111146 705242 111382 705478
rect 110826 669218 111062 669454
rect 111146 669218 111382 669454
rect 110826 668898 111062 669134
rect 111146 668898 111382 669134
rect 110826 633218 111062 633454
rect 111146 633218 111382 633454
rect 110826 632898 111062 633134
rect 111146 632898 111382 633134
rect 110826 597218 111062 597454
rect 111146 597218 111382 597454
rect 110826 596898 111062 597134
rect 111146 596898 111382 597134
rect 110826 561218 111062 561454
rect 111146 561218 111382 561454
rect 110826 560898 111062 561134
rect 111146 560898 111382 561134
rect 110826 525218 111062 525454
rect 111146 525218 111382 525454
rect 110826 524898 111062 525134
rect 111146 524898 111382 525134
rect 110826 489218 111062 489454
rect 111146 489218 111382 489454
rect 110826 488898 111062 489134
rect 111146 488898 111382 489134
rect 110826 453218 111062 453454
rect 111146 453218 111382 453454
rect 110826 452898 111062 453134
rect 111146 452898 111382 453134
rect 110826 417218 111062 417454
rect 111146 417218 111382 417454
rect 110826 416898 111062 417134
rect 111146 416898 111382 417134
rect 110826 381218 111062 381454
rect 111146 381218 111382 381454
rect 110826 380898 111062 381134
rect 111146 380898 111382 381134
rect 110826 345218 111062 345454
rect 111146 345218 111382 345454
rect 110826 344898 111062 345134
rect 111146 344898 111382 345134
rect 110826 309218 111062 309454
rect 111146 309218 111382 309454
rect 110826 308898 111062 309134
rect 111146 308898 111382 309134
rect 110826 273218 111062 273454
rect 111146 273218 111382 273454
rect 110826 272898 111062 273134
rect 111146 272898 111382 273134
rect 110826 237218 111062 237454
rect 111146 237218 111382 237454
rect 110826 236898 111062 237134
rect 111146 236898 111382 237134
rect 110826 201218 111062 201454
rect 111146 201218 111382 201454
rect 110826 200898 111062 201134
rect 111146 200898 111382 201134
rect 110826 165218 111062 165454
rect 111146 165218 111382 165454
rect 110826 164898 111062 165134
rect 111146 164898 111382 165134
rect 110826 129218 111062 129454
rect 111146 129218 111382 129454
rect 110826 128898 111062 129134
rect 111146 128898 111382 129134
rect 110826 93218 111062 93454
rect 111146 93218 111382 93454
rect 110826 92898 111062 93134
rect 111146 92898 111382 93134
rect 110826 57218 111062 57454
rect 111146 57218 111382 57454
rect 110826 56898 111062 57134
rect 111146 56898 111382 57134
rect 110826 21218 111062 21454
rect 111146 21218 111382 21454
rect 110826 20898 111062 21134
rect 111146 20898 111382 21134
rect 110826 -1542 111062 -1306
rect 111146 -1542 111382 -1306
rect 110826 -1862 111062 -1626
rect 111146 -1862 111382 -1626
rect 121986 711322 122222 711558
rect 122306 711322 122542 711558
rect 121986 711002 122222 711238
rect 122306 711002 122542 711238
rect 118266 709402 118502 709638
rect 118586 709402 118822 709638
rect 118266 709082 118502 709318
rect 118586 709082 118822 709318
rect 111986 698378 112222 698614
rect 112306 698378 112542 698614
rect 111986 698058 112222 698294
rect 112306 698058 112542 698294
rect 111986 662378 112222 662614
rect 112306 662378 112542 662614
rect 111986 662058 112222 662294
rect 112306 662058 112542 662294
rect 111986 626378 112222 626614
rect 112306 626378 112542 626614
rect 111986 626058 112222 626294
rect 112306 626058 112542 626294
rect 111986 590378 112222 590614
rect 112306 590378 112542 590614
rect 111986 590058 112222 590294
rect 112306 590058 112542 590294
rect 111986 554378 112222 554614
rect 112306 554378 112542 554614
rect 111986 554058 112222 554294
rect 112306 554058 112542 554294
rect 111986 518378 112222 518614
rect 112306 518378 112542 518614
rect 111986 518058 112222 518294
rect 112306 518058 112542 518294
rect 111986 482378 112222 482614
rect 112306 482378 112542 482614
rect 111986 482058 112222 482294
rect 112306 482058 112542 482294
rect 111986 446378 112222 446614
rect 112306 446378 112542 446614
rect 111986 446058 112222 446294
rect 112306 446058 112542 446294
rect 111986 410378 112222 410614
rect 112306 410378 112542 410614
rect 111986 410058 112222 410294
rect 112306 410058 112542 410294
rect 111986 374378 112222 374614
rect 112306 374378 112542 374614
rect 111986 374058 112222 374294
rect 112306 374058 112542 374294
rect 111986 338378 112222 338614
rect 112306 338378 112542 338614
rect 111986 338058 112222 338294
rect 112306 338058 112542 338294
rect 111986 302378 112222 302614
rect 112306 302378 112542 302614
rect 111986 302058 112222 302294
rect 112306 302058 112542 302294
rect 111986 266378 112222 266614
rect 112306 266378 112542 266614
rect 111986 266058 112222 266294
rect 112306 266058 112542 266294
rect 111986 230378 112222 230614
rect 112306 230378 112542 230614
rect 111986 230058 112222 230294
rect 112306 230058 112542 230294
rect 111986 194378 112222 194614
rect 112306 194378 112542 194614
rect 111986 194058 112222 194294
rect 112306 194058 112542 194294
rect 111986 158378 112222 158614
rect 112306 158378 112542 158614
rect 111986 158058 112222 158294
rect 112306 158058 112542 158294
rect 111986 122378 112222 122614
rect 112306 122378 112542 122614
rect 111986 122058 112222 122294
rect 112306 122058 112542 122294
rect 111986 86378 112222 86614
rect 112306 86378 112542 86614
rect 111986 86058 112222 86294
rect 112306 86058 112542 86294
rect 111986 50378 112222 50614
rect 112306 50378 112542 50614
rect 111986 50058 112222 50294
rect 112306 50058 112542 50294
rect 111986 14378 112222 14614
rect 112306 14378 112542 14614
rect 111986 14058 112222 14294
rect 112306 14058 112542 14294
rect 108266 -4422 108502 -4186
rect 108586 -4422 108822 -4186
rect 108266 -4742 108502 -4506
rect 108586 -4742 108822 -4506
rect 101986 -7302 102222 -7066
rect 102306 -7302 102542 -7066
rect 101986 -7622 102222 -7386
rect 102306 -7622 102542 -7386
rect 114546 707482 114782 707718
rect 114866 707482 115102 707718
rect 114546 707162 114782 707398
rect 114866 707162 115102 707398
rect 114546 672938 114782 673174
rect 114866 672938 115102 673174
rect 114546 672618 114782 672854
rect 114866 672618 115102 672854
rect 114546 636938 114782 637174
rect 114866 636938 115102 637174
rect 114546 636618 114782 636854
rect 114866 636618 115102 636854
rect 114546 600938 114782 601174
rect 114866 600938 115102 601174
rect 114546 600618 114782 600854
rect 114866 600618 115102 600854
rect 114546 564938 114782 565174
rect 114866 564938 115102 565174
rect 114546 564618 114782 564854
rect 114866 564618 115102 564854
rect 114546 528938 114782 529174
rect 114866 528938 115102 529174
rect 114546 528618 114782 528854
rect 114866 528618 115102 528854
rect 114546 492938 114782 493174
rect 114866 492938 115102 493174
rect 114546 492618 114782 492854
rect 114866 492618 115102 492854
rect 114546 456938 114782 457174
rect 114866 456938 115102 457174
rect 114546 456618 114782 456854
rect 114866 456618 115102 456854
rect 114546 420938 114782 421174
rect 114866 420938 115102 421174
rect 114546 420618 114782 420854
rect 114866 420618 115102 420854
rect 114546 384938 114782 385174
rect 114866 384938 115102 385174
rect 114546 384618 114782 384854
rect 114866 384618 115102 384854
rect 114546 348938 114782 349174
rect 114866 348938 115102 349174
rect 114546 348618 114782 348854
rect 114866 348618 115102 348854
rect 114546 312938 114782 313174
rect 114866 312938 115102 313174
rect 114546 312618 114782 312854
rect 114866 312618 115102 312854
rect 114546 276938 114782 277174
rect 114866 276938 115102 277174
rect 114546 276618 114782 276854
rect 114866 276618 115102 276854
rect 114546 240938 114782 241174
rect 114866 240938 115102 241174
rect 114546 240618 114782 240854
rect 114866 240618 115102 240854
rect 114546 204938 114782 205174
rect 114866 204938 115102 205174
rect 114546 204618 114782 204854
rect 114866 204618 115102 204854
rect 114546 168938 114782 169174
rect 114866 168938 115102 169174
rect 114546 168618 114782 168854
rect 114866 168618 115102 168854
rect 114546 132938 114782 133174
rect 114866 132938 115102 133174
rect 114546 132618 114782 132854
rect 114866 132618 115102 132854
rect 114546 96938 114782 97174
rect 114866 96938 115102 97174
rect 114546 96618 114782 96854
rect 114866 96618 115102 96854
rect 114546 60938 114782 61174
rect 114866 60938 115102 61174
rect 114546 60618 114782 60854
rect 114866 60618 115102 60854
rect 114546 24938 114782 25174
rect 114866 24938 115102 25174
rect 114546 24618 114782 24854
rect 114866 24618 115102 24854
rect 114546 -3462 114782 -3226
rect 114866 -3462 115102 -3226
rect 114546 -3782 114782 -3546
rect 114866 -3782 115102 -3546
rect 118266 676658 118502 676894
rect 118586 676658 118822 676894
rect 118266 676338 118502 676574
rect 118586 676338 118822 676574
rect 118266 640658 118502 640894
rect 118586 640658 118822 640894
rect 118266 640338 118502 640574
rect 118586 640338 118822 640574
rect 118266 604658 118502 604894
rect 118586 604658 118822 604894
rect 118266 604338 118502 604574
rect 118586 604338 118822 604574
rect 118266 568658 118502 568894
rect 118586 568658 118822 568894
rect 118266 568338 118502 568574
rect 118586 568338 118822 568574
rect 118266 532658 118502 532894
rect 118586 532658 118822 532894
rect 118266 532338 118502 532574
rect 118586 532338 118822 532574
rect 118266 496658 118502 496894
rect 118586 496658 118822 496894
rect 118266 496338 118502 496574
rect 118586 496338 118822 496574
rect 118266 460658 118502 460894
rect 118586 460658 118822 460894
rect 118266 460338 118502 460574
rect 118586 460338 118822 460574
rect 118266 424658 118502 424894
rect 118586 424658 118822 424894
rect 118266 424338 118502 424574
rect 118586 424338 118822 424574
rect 118266 388658 118502 388894
rect 118586 388658 118822 388894
rect 118266 388338 118502 388574
rect 118586 388338 118822 388574
rect 118266 352658 118502 352894
rect 118586 352658 118822 352894
rect 118266 352338 118502 352574
rect 118586 352338 118822 352574
rect 118266 316658 118502 316894
rect 118586 316658 118822 316894
rect 118266 316338 118502 316574
rect 118586 316338 118822 316574
rect 118266 280658 118502 280894
rect 118586 280658 118822 280894
rect 118266 280338 118502 280574
rect 118586 280338 118822 280574
rect 118266 244658 118502 244894
rect 118586 244658 118822 244894
rect 118266 244338 118502 244574
rect 118586 244338 118822 244574
rect 118266 208658 118502 208894
rect 118586 208658 118822 208894
rect 118266 208338 118502 208574
rect 118586 208338 118822 208574
rect 118266 172658 118502 172894
rect 118586 172658 118822 172894
rect 118266 172338 118502 172574
rect 118586 172338 118822 172574
rect 118266 136658 118502 136894
rect 118586 136658 118822 136894
rect 118266 136338 118502 136574
rect 118586 136338 118822 136574
rect 118266 100658 118502 100894
rect 118586 100658 118822 100894
rect 118266 100338 118502 100574
rect 118586 100338 118822 100574
rect 118266 64658 118502 64894
rect 118586 64658 118822 64894
rect 118266 64338 118502 64574
rect 118586 64338 118822 64574
rect 118266 28658 118502 28894
rect 118586 28658 118822 28894
rect 118266 28338 118502 28574
rect 118586 28338 118822 28574
rect 120826 704602 121062 704838
rect 121146 704602 121382 704838
rect 120826 704282 121062 704518
rect 121146 704282 121382 704518
rect 120826 687218 121062 687454
rect 121146 687218 121382 687454
rect 120826 686898 121062 687134
rect 121146 686898 121382 687134
rect 120826 651218 121062 651454
rect 121146 651218 121382 651454
rect 120826 650898 121062 651134
rect 121146 650898 121382 651134
rect 120826 615218 121062 615454
rect 121146 615218 121382 615454
rect 120826 614898 121062 615134
rect 121146 614898 121382 615134
rect 120826 579218 121062 579454
rect 121146 579218 121382 579454
rect 120826 578898 121062 579134
rect 121146 578898 121382 579134
rect 120826 543218 121062 543454
rect 121146 543218 121382 543454
rect 120826 542898 121062 543134
rect 121146 542898 121382 543134
rect 120826 507218 121062 507454
rect 121146 507218 121382 507454
rect 120826 506898 121062 507134
rect 121146 506898 121382 507134
rect 120826 471218 121062 471454
rect 121146 471218 121382 471454
rect 120826 470898 121062 471134
rect 121146 470898 121382 471134
rect 120826 435218 121062 435454
rect 121146 435218 121382 435454
rect 120826 434898 121062 435134
rect 121146 434898 121382 435134
rect 120826 399218 121062 399454
rect 121146 399218 121382 399454
rect 120826 398898 121062 399134
rect 121146 398898 121382 399134
rect 120826 363218 121062 363454
rect 121146 363218 121382 363454
rect 120826 362898 121062 363134
rect 121146 362898 121382 363134
rect 120826 327218 121062 327454
rect 121146 327218 121382 327454
rect 120826 326898 121062 327134
rect 121146 326898 121382 327134
rect 120826 291218 121062 291454
rect 121146 291218 121382 291454
rect 120826 290898 121062 291134
rect 121146 290898 121382 291134
rect 120826 255218 121062 255454
rect 121146 255218 121382 255454
rect 120826 254898 121062 255134
rect 121146 254898 121382 255134
rect 120826 219218 121062 219454
rect 121146 219218 121382 219454
rect 120826 218898 121062 219134
rect 121146 218898 121382 219134
rect 120826 183218 121062 183454
rect 121146 183218 121382 183454
rect 120826 182898 121062 183134
rect 121146 182898 121382 183134
rect 120826 147218 121062 147454
rect 121146 147218 121382 147454
rect 120826 146898 121062 147134
rect 121146 146898 121382 147134
rect 120826 111218 121062 111454
rect 121146 111218 121382 111454
rect 120826 110898 121062 111134
rect 121146 110898 121382 111134
rect 120826 75218 121062 75454
rect 121146 75218 121382 75454
rect 120826 74898 121062 75134
rect 121146 74898 121382 75134
rect 120826 39218 121062 39454
rect 121146 39218 121382 39454
rect 120826 38898 121062 39134
rect 121146 38898 121382 39134
rect 120826 3218 121062 3454
rect 121146 3218 121382 3454
rect 120826 2898 121062 3134
rect 121146 2898 121382 3134
rect 120826 -582 121062 -346
rect 121146 -582 121382 -346
rect 120826 -902 121062 -666
rect 121146 -902 121382 -666
rect 131986 710362 132222 710598
rect 132306 710362 132542 710598
rect 131986 710042 132222 710278
rect 132306 710042 132542 710278
rect 128266 708442 128502 708678
rect 128586 708442 128822 708678
rect 128266 708122 128502 708358
rect 128586 708122 128822 708358
rect 121986 680378 122222 680614
rect 122306 680378 122542 680614
rect 121986 680058 122222 680294
rect 122306 680058 122542 680294
rect 121986 644378 122222 644614
rect 122306 644378 122542 644614
rect 121986 644058 122222 644294
rect 122306 644058 122542 644294
rect 121986 608378 122222 608614
rect 122306 608378 122542 608614
rect 121986 608058 122222 608294
rect 122306 608058 122542 608294
rect 121986 572378 122222 572614
rect 122306 572378 122542 572614
rect 121986 572058 122222 572294
rect 122306 572058 122542 572294
rect 121986 536378 122222 536614
rect 122306 536378 122542 536614
rect 121986 536058 122222 536294
rect 122306 536058 122542 536294
rect 121986 500378 122222 500614
rect 122306 500378 122542 500614
rect 121986 500058 122222 500294
rect 122306 500058 122542 500294
rect 121986 464378 122222 464614
rect 122306 464378 122542 464614
rect 121986 464058 122222 464294
rect 122306 464058 122542 464294
rect 121986 428378 122222 428614
rect 122306 428378 122542 428614
rect 121986 428058 122222 428294
rect 122306 428058 122542 428294
rect 121986 392378 122222 392614
rect 122306 392378 122542 392614
rect 121986 392058 122222 392294
rect 122306 392058 122542 392294
rect 121986 356378 122222 356614
rect 122306 356378 122542 356614
rect 121986 356058 122222 356294
rect 122306 356058 122542 356294
rect 121986 320378 122222 320614
rect 122306 320378 122542 320614
rect 121986 320058 122222 320294
rect 122306 320058 122542 320294
rect 121986 284378 122222 284614
rect 122306 284378 122542 284614
rect 121986 284058 122222 284294
rect 122306 284058 122542 284294
rect 121986 248378 122222 248614
rect 122306 248378 122542 248614
rect 121986 248058 122222 248294
rect 122306 248058 122542 248294
rect 121986 212378 122222 212614
rect 122306 212378 122542 212614
rect 121986 212058 122222 212294
rect 122306 212058 122542 212294
rect 121986 176378 122222 176614
rect 122306 176378 122542 176614
rect 121986 176058 122222 176294
rect 122306 176058 122542 176294
rect 121986 140378 122222 140614
rect 122306 140378 122542 140614
rect 121986 140058 122222 140294
rect 122306 140058 122542 140294
rect 121986 104378 122222 104614
rect 122306 104378 122542 104614
rect 121986 104058 122222 104294
rect 122306 104058 122542 104294
rect 121986 68378 122222 68614
rect 122306 68378 122542 68614
rect 121986 68058 122222 68294
rect 122306 68058 122542 68294
rect 121986 32378 122222 32614
rect 122306 32378 122542 32614
rect 121986 32058 122222 32294
rect 122306 32058 122542 32294
rect 118266 -5382 118502 -5146
rect 118586 -5382 118822 -5146
rect 118266 -5702 118502 -5466
rect 118586 -5702 118822 -5466
rect 111986 -6342 112222 -6106
rect 112306 -6342 112542 -6106
rect 111986 -6662 112222 -6426
rect 112306 -6662 112542 -6426
rect 124546 706522 124782 706758
rect 124866 706522 125102 706758
rect 124546 706202 124782 706438
rect 124866 706202 125102 706438
rect 124546 690938 124782 691174
rect 124866 690938 125102 691174
rect 124546 690618 124782 690854
rect 124866 690618 125102 690854
rect 124546 654938 124782 655174
rect 124866 654938 125102 655174
rect 124546 654618 124782 654854
rect 124866 654618 125102 654854
rect 124546 618938 124782 619174
rect 124866 618938 125102 619174
rect 124546 618618 124782 618854
rect 124866 618618 125102 618854
rect 124546 582938 124782 583174
rect 124866 582938 125102 583174
rect 124546 582618 124782 582854
rect 124866 582618 125102 582854
rect 124546 546938 124782 547174
rect 124866 546938 125102 547174
rect 124546 546618 124782 546854
rect 124866 546618 125102 546854
rect 124546 510938 124782 511174
rect 124866 510938 125102 511174
rect 124546 510618 124782 510854
rect 124866 510618 125102 510854
rect 124546 474938 124782 475174
rect 124866 474938 125102 475174
rect 124546 474618 124782 474854
rect 124866 474618 125102 474854
rect 124546 438938 124782 439174
rect 124866 438938 125102 439174
rect 124546 438618 124782 438854
rect 124866 438618 125102 438854
rect 124546 402938 124782 403174
rect 124866 402938 125102 403174
rect 124546 402618 124782 402854
rect 124866 402618 125102 402854
rect 124546 366938 124782 367174
rect 124866 366938 125102 367174
rect 124546 366618 124782 366854
rect 124866 366618 125102 366854
rect 124546 330938 124782 331174
rect 124866 330938 125102 331174
rect 124546 330618 124782 330854
rect 124866 330618 125102 330854
rect 124546 294938 124782 295174
rect 124866 294938 125102 295174
rect 124546 294618 124782 294854
rect 124866 294618 125102 294854
rect 124546 258938 124782 259174
rect 124866 258938 125102 259174
rect 124546 258618 124782 258854
rect 124866 258618 125102 258854
rect 124546 222938 124782 223174
rect 124866 222938 125102 223174
rect 124546 222618 124782 222854
rect 124866 222618 125102 222854
rect 124546 186938 124782 187174
rect 124866 186938 125102 187174
rect 124546 186618 124782 186854
rect 124866 186618 125102 186854
rect 124546 150938 124782 151174
rect 124866 150938 125102 151174
rect 124546 150618 124782 150854
rect 124866 150618 125102 150854
rect 124546 114938 124782 115174
rect 124866 114938 125102 115174
rect 124546 114618 124782 114854
rect 124866 114618 125102 114854
rect 124546 78938 124782 79174
rect 124866 78938 125102 79174
rect 124546 78618 124782 78854
rect 124866 78618 125102 78854
rect 124546 42938 124782 43174
rect 124866 42938 125102 43174
rect 124546 42618 124782 42854
rect 124866 42618 125102 42854
rect 124546 6938 124782 7174
rect 124866 6938 125102 7174
rect 124546 6618 124782 6854
rect 124866 6618 125102 6854
rect 124546 -2502 124782 -2266
rect 124866 -2502 125102 -2266
rect 124546 -2822 124782 -2586
rect 124866 -2822 125102 -2586
rect 128266 694658 128502 694894
rect 128586 694658 128822 694894
rect 128266 694338 128502 694574
rect 128586 694338 128822 694574
rect 128266 658658 128502 658894
rect 128586 658658 128822 658894
rect 128266 658338 128502 658574
rect 128586 658338 128822 658574
rect 128266 622658 128502 622894
rect 128586 622658 128822 622894
rect 128266 622338 128502 622574
rect 128586 622338 128822 622574
rect 128266 586658 128502 586894
rect 128586 586658 128822 586894
rect 128266 586338 128502 586574
rect 128586 586338 128822 586574
rect 128266 550658 128502 550894
rect 128586 550658 128822 550894
rect 128266 550338 128502 550574
rect 128586 550338 128822 550574
rect 128266 514658 128502 514894
rect 128586 514658 128822 514894
rect 128266 514338 128502 514574
rect 128586 514338 128822 514574
rect 128266 478658 128502 478894
rect 128586 478658 128822 478894
rect 128266 478338 128502 478574
rect 128586 478338 128822 478574
rect 128266 442658 128502 442894
rect 128586 442658 128822 442894
rect 128266 442338 128502 442574
rect 128586 442338 128822 442574
rect 128266 406658 128502 406894
rect 128586 406658 128822 406894
rect 128266 406338 128502 406574
rect 128586 406338 128822 406574
rect 128266 370658 128502 370894
rect 128586 370658 128822 370894
rect 128266 370338 128502 370574
rect 128586 370338 128822 370574
rect 128266 334658 128502 334894
rect 128586 334658 128822 334894
rect 128266 334338 128502 334574
rect 128586 334338 128822 334574
rect 128266 298658 128502 298894
rect 128586 298658 128822 298894
rect 128266 298338 128502 298574
rect 128586 298338 128822 298574
rect 128266 262658 128502 262894
rect 128586 262658 128822 262894
rect 128266 262338 128502 262574
rect 128586 262338 128822 262574
rect 128266 226658 128502 226894
rect 128586 226658 128822 226894
rect 128266 226338 128502 226574
rect 128586 226338 128822 226574
rect 128266 190658 128502 190894
rect 128586 190658 128822 190894
rect 128266 190338 128502 190574
rect 128586 190338 128822 190574
rect 128266 154658 128502 154894
rect 128586 154658 128822 154894
rect 128266 154338 128502 154574
rect 128586 154338 128822 154574
rect 128266 118658 128502 118894
rect 128586 118658 128822 118894
rect 128266 118338 128502 118574
rect 128586 118338 128822 118574
rect 128266 82658 128502 82894
rect 128586 82658 128822 82894
rect 128266 82338 128502 82574
rect 128586 82338 128822 82574
rect 128266 46658 128502 46894
rect 128586 46658 128822 46894
rect 128266 46338 128502 46574
rect 128586 46338 128822 46574
rect 128266 10658 128502 10894
rect 128586 10658 128822 10894
rect 128266 10338 128502 10574
rect 128586 10338 128822 10574
rect 130826 705562 131062 705798
rect 131146 705562 131382 705798
rect 130826 705242 131062 705478
rect 131146 705242 131382 705478
rect 130826 669218 131062 669454
rect 131146 669218 131382 669454
rect 130826 668898 131062 669134
rect 131146 668898 131382 669134
rect 130826 633218 131062 633454
rect 131146 633218 131382 633454
rect 130826 632898 131062 633134
rect 131146 632898 131382 633134
rect 130826 597218 131062 597454
rect 131146 597218 131382 597454
rect 130826 596898 131062 597134
rect 131146 596898 131382 597134
rect 130826 561218 131062 561454
rect 131146 561218 131382 561454
rect 130826 560898 131062 561134
rect 131146 560898 131382 561134
rect 130826 525218 131062 525454
rect 131146 525218 131382 525454
rect 130826 524898 131062 525134
rect 131146 524898 131382 525134
rect 130826 489218 131062 489454
rect 131146 489218 131382 489454
rect 130826 488898 131062 489134
rect 131146 488898 131382 489134
rect 130826 453218 131062 453454
rect 131146 453218 131382 453454
rect 130826 452898 131062 453134
rect 131146 452898 131382 453134
rect 130826 417218 131062 417454
rect 131146 417218 131382 417454
rect 130826 416898 131062 417134
rect 131146 416898 131382 417134
rect 130826 381218 131062 381454
rect 131146 381218 131382 381454
rect 130826 380898 131062 381134
rect 131146 380898 131382 381134
rect 130826 345218 131062 345454
rect 131146 345218 131382 345454
rect 130826 344898 131062 345134
rect 131146 344898 131382 345134
rect 130826 309218 131062 309454
rect 131146 309218 131382 309454
rect 130826 308898 131062 309134
rect 131146 308898 131382 309134
rect 130826 273218 131062 273454
rect 131146 273218 131382 273454
rect 130826 272898 131062 273134
rect 131146 272898 131382 273134
rect 130826 237218 131062 237454
rect 131146 237218 131382 237454
rect 130826 236898 131062 237134
rect 131146 236898 131382 237134
rect 130826 201218 131062 201454
rect 131146 201218 131382 201454
rect 130826 200898 131062 201134
rect 131146 200898 131382 201134
rect 130826 165218 131062 165454
rect 131146 165218 131382 165454
rect 130826 164898 131062 165134
rect 131146 164898 131382 165134
rect 130826 129218 131062 129454
rect 131146 129218 131382 129454
rect 130826 128898 131062 129134
rect 131146 128898 131382 129134
rect 130826 93218 131062 93454
rect 131146 93218 131382 93454
rect 130826 92898 131062 93134
rect 131146 92898 131382 93134
rect 130826 57218 131062 57454
rect 131146 57218 131382 57454
rect 130826 56898 131062 57134
rect 131146 56898 131382 57134
rect 130826 21218 131062 21454
rect 131146 21218 131382 21454
rect 130826 20898 131062 21134
rect 131146 20898 131382 21134
rect 130826 -1542 131062 -1306
rect 131146 -1542 131382 -1306
rect 130826 -1862 131062 -1626
rect 131146 -1862 131382 -1626
rect 141986 711322 142222 711558
rect 142306 711322 142542 711558
rect 141986 711002 142222 711238
rect 142306 711002 142542 711238
rect 138266 709402 138502 709638
rect 138586 709402 138822 709638
rect 138266 709082 138502 709318
rect 138586 709082 138822 709318
rect 131986 698378 132222 698614
rect 132306 698378 132542 698614
rect 131986 698058 132222 698294
rect 132306 698058 132542 698294
rect 131986 662378 132222 662614
rect 132306 662378 132542 662614
rect 131986 662058 132222 662294
rect 132306 662058 132542 662294
rect 131986 626378 132222 626614
rect 132306 626378 132542 626614
rect 131986 626058 132222 626294
rect 132306 626058 132542 626294
rect 131986 590378 132222 590614
rect 132306 590378 132542 590614
rect 131986 590058 132222 590294
rect 132306 590058 132542 590294
rect 131986 554378 132222 554614
rect 132306 554378 132542 554614
rect 131986 554058 132222 554294
rect 132306 554058 132542 554294
rect 131986 518378 132222 518614
rect 132306 518378 132542 518614
rect 131986 518058 132222 518294
rect 132306 518058 132542 518294
rect 131986 482378 132222 482614
rect 132306 482378 132542 482614
rect 131986 482058 132222 482294
rect 132306 482058 132542 482294
rect 131986 446378 132222 446614
rect 132306 446378 132542 446614
rect 131986 446058 132222 446294
rect 132306 446058 132542 446294
rect 131986 410378 132222 410614
rect 132306 410378 132542 410614
rect 131986 410058 132222 410294
rect 132306 410058 132542 410294
rect 131986 374378 132222 374614
rect 132306 374378 132542 374614
rect 131986 374058 132222 374294
rect 132306 374058 132542 374294
rect 131986 338378 132222 338614
rect 132306 338378 132542 338614
rect 131986 338058 132222 338294
rect 132306 338058 132542 338294
rect 131986 302378 132222 302614
rect 132306 302378 132542 302614
rect 131986 302058 132222 302294
rect 132306 302058 132542 302294
rect 131986 266378 132222 266614
rect 132306 266378 132542 266614
rect 131986 266058 132222 266294
rect 132306 266058 132542 266294
rect 131986 230378 132222 230614
rect 132306 230378 132542 230614
rect 131986 230058 132222 230294
rect 132306 230058 132542 230294
rect 131986 194378 132222 194614
rect 132306 194378 132542 194614
rect 131986 194058 132222 194294
rect 132306 194058 132542 194294
rect 131986 158378 132222 158614
rect 132306 158378 132542 158614
rect 131986 158058 132222 158294
rect 132306 158058 132542 158294
rect 131986 122378 132222 122614
rect 132306 122378 132542 122614
rect 131986 122058 132222 122294
rect 132306 122058 132542 122294
rect 131986 86378 132222 86614
rect 132306 86378 132542 86614
rect 131986 86058 132222 86294
rect 132306 86058 132542 86294
rect 131986 50378 132222 50614
rect 132306 50378 132542 50614
rect 131986 50058 132222 50294
rect 132306 50058 132542 50294
rect 131986 14378 132222 14614
rect 132306 14378 132542 14614
rect 131986 14058 132222 14294
rect 132306 14058 132542 14294
rect 128266 -4422 128502 -4186
rect 128586 -4422 128822 -4186
rect 128266 -4742 128502 -4506
rect 128586 -4742 128822 -4506
rect 121986 -7302 122222 -7066
rect 122306 -7302 122542 -7066
rect 121986 -7622 122222 -7386
rect 122306 -7622 122542 -7386
rect 134546 707482 134782 707718
rect 134866 707482 135102 707718
rect 134546 707162 134782 707398
rect 134866 707162 135102 707398
rect 134546 672938 134782 673174
rect 134866 672938 135102 673174
rect 134546 672618 134782 672854
rect 134866 672618 135102 672854
rect 134546 636938 134782 637174
rect 134866 636938 135102 637174
rect 134546 636618 134782 636854
rect 134866 636618 135102 636854
rect 134546 600938 134782 601174
rect 134866 600938 135102 601174
rect 134546 600618 134782 600854
rect 134866 600618 135102 600854
rect 134546 564938 134782 565174
rect 134866 564938 135102 565174
rect 134546 564618 134782 564854
rect 134866 564618 135102 564854
rect 134546 528938 134782 529174
rect 134866 528938 135102 529174
rect 134546 528618 134782 528854
rect 134866 528618 135102 528854
rect 134546 492938 134782 493174
rect 134866 492938 135102 493174
rect 134546 492618 134782 492854
rect 134866 492618 135102 492854
rect 134546 456938 134782 457174
rect 134866 456938 135102 457174
rect 134546 456618 134782 456854
rect 134866 456618 135102 456854
rect 134546 420938 134782 421174
rect 134866 420938 135102 421174
rect 134546 420618 134782 420854
rect 134866 420618 135102 420854
rect 134546 384938 134782 385174
rect 134866 384938 135102 385174
rect 134546 384618 134782 384854
rect 134866 384618 135102 384854
rect 134546 348938 134782 349174
rect 134866 348938 135102 349174
rect 134546 348618 134782 348854
rect 134866 348618 135102 348854
rect 134546 312938 134782 313174
rect 134866 312938 135102 313174
rect 134546 312618 134782 312854
rect 134866 312618 135102 312854
rect 134546 276938 134782 277174
rect 134866 276938 135102 277174
rect 134546 276618 134782 276854
rect 134866 276618 135102 276854
rect 134546 240938 134782 241174
rect 134866 240938 135102 241174
rect 134546 240618 134782 240854
rect 134866 240618 135102 240854
rect 134546 204938 134782 205174
rect 134866 204938 135102 205174
rect 134546 204618 134782 204854
rect 134866 204618 135102 204854
rect 134546 168938 134782 169174
rect 134866 168938 135102 169174
rect 134546 168618 134782 168854
rect 134866 168618 135102 168854
rect 134546 132938 134782 133174
rect 134866 132938 135102 133174
rect 134546 132618 134782 132854
rect 134866 132618 135102 132854
rect 134546 96938 134782 97174
rect 134866 96938 135102 97174
rect 134546 96618 134782 96854
rect 134866 96618 135102 96854
rect 134546 60938 134782 61174
rect 134866 60938 135102 61174
rect 134546 60618 134782 60854
rect 134866 60618 135102 60854
rect 134546 24938 134782 25174
rect 134866 24938 135102 25174
rect 134546 24618 134782 24854
rect 134866 24618 135102 24854
rect 134546 -3462 134782 -3226
rect 134866 -3462 135102 -3226
rect 134546 -3782 134782 -3546
rect 134866 -3782 135102 -3546
rect 138266 676658 138502 676894
rect 138586 676658 138822 676894
rect 138266 676338 138502 676574
rect 138586 676338 138822 676574
rect 138266 640658 138502 640894
rect 138586 640658 138822 640894
rect 138266 640338 138502 640574
rect 138586 640338 138822 640574
rect 138266 604658 138502 604894
rect 138586 604658 138822 604894
rect 138266 604338 138502 604574
rect 138586 604338 138822 604574
rect 138266 568658 138502 568894
rect 138586 568658 138822 568894
rect 138266 568338 138502 568574
rect 138586 568338 138822 568574
rect 138266 532658 138502 532894
rect 138586 532658 138822 532894
rect 138266 532338 138502 532574
rect 138586 532338 138822 532574
rect 138266 496658 138502 496894
rect 138586 496658 138822 496894
rect 138266 496338 138502 496574
rect 138586 496338 138822 496574
rect 138266 460658 138502 460894
rect 138586 460658 138822 460894
rect 138266 460338 138502 460574
rect 138586 460338 138822 460574
rect 138266 424658 138502 424894
rect 138586 424658 138822 424894
rect 138266 424338 138502 424574
rect 138586 424338 138822 424574
rect 138266 388658 138502 388894
rect 138586 388658 138822 388894
rect 138266 388338 138502 388574
rect 138586 388338 138822 388574
rect 138266 352658 138502 352894
rect 138586 352658 138822 352894
rect 138266 352338 138502 352574
rect 138586 352338 138822 352574
rect 138266 316658 138502 316894
rect 138586 316658 138822 316894
rect 138266 316338 138502 316574
rect 138586 316338 138822 316574
rect 138266 280658 138502 280894
rect 138586 280658 138822 280894
rect 138266 280338 138502 280574
rect 138586 280338 138822 280574
rect 138266 244658 138502 244894
rect 138586 244658 138822 244894
rect 138266 244338 138502 244574
rect 138586 244338 138822 244574
rect 138266 208658 138502 208894
rect 138586 208658 138822 208894
rect 138266 208338 138502 208574
rect 138586 208338 138822 208574
rect 138266 172658 138502 172894
rect 138586 172658 138822 172894
rect 138266 172338 138502 172574
rect 138586 172338 138822 172574
rect 138266 136658 138502 136894
rect 138586 136658 138822 136894
rect 138266 136338 138502 136574
rect 138586 136338 138822 136574
rect 138266 100658 138502 100894
rect 138586 100658 138822 100894
rect 138266 100338 138502 100574
rect 138586 100338 138822 100574
rect 138266 64658 138502 64894
rect 138586 64658 138822 64894
rect 138266 64338 138502 64574
rect 138586 64338 138822 64574
rect 138266 28658 138502 28894
rect 138586 28658 138822 28894
rect 138266 28338 138502 28574
rect 138586 28338 138822 28574
rect 140826 704602 141062 704838
rect 141146 704602 141382 704838
rect 140826 704282 141062 704518
rect 141146 704282 141382 704518
rect 140826 687218 141062 687454
rect 141146 687218 141382 687454
rect 140826 686898 141062 687134
rect 141146 686898 141382 687134
rect 140826 651218 141062 651454
rect 141146 651218 141382 651454
rect 140826 650898 141062 651134
rect 141146 650898 141382 651134
rect 140826 615218 141062 615454
rect 141146 615218 141382 615454
rect 140826 614898 141062 615134
rect 141146 614898 141382 615134
rect 140826 579218 141062 579454
rect 141146 579218 141382 579454
rect 140826 578898 141062 579134
rect 141146 578898 141382 579134
rect 140826 543218 141062 543454
rect 141146 543218 141382 543454
rect 140826 542898 141062 543134
rect 141146 542898 141382 543134
rect 140826 507218 141062 507454
rect 141146 507218 141382 507454
rect 140826 506898 141062 507134
rect 141146 506898 141382 507134
rect 140826 471218 141062 471454
rect 141146 471218 141382 471454
rect 140826 470898 141062 471134
rect 141146 470898 141382 471134
rect 140826 435218 141062 435454
rect 141146 435218 141382 435454
rect 140826 434898 141062 435134
rect 141146 434898 141382 435134
rect 140826 399218 141062 399454
rect 141146 399218 141382 399454
rect 140826 398898 141062 399134
rect 141146 398898 141382 399134
rect 140826 363218 141062 363454
rect 141146 363218 141382 363454
rect 140826 362898 141062 363134
rect 141146 362898 141382 363134
rect 140826 327218 141062 327454
rect 141146 327218 141382 327454
rect 140826 326898 141062 327134
rect 141146 326898 141382 327134
rect 140826 291218 141062 291454
rect 141146 291218 141382 291454
rect 140826 290898 141062 291134
rect 141146 290898 141382 291134
rect 140826 255218 141062 255454
rect 141146 255218 141382 255454
rect 140826 254898 141062 255134
rect 141146 254898 141382 255134
rect 140826 219218 141062 219454
rect 141146 219218 141382 219454
rect 140826 218898 141062 219134
rect 141146 218898 141382 219134
rect 140826 183218 141062 183454
rect 141146 183218 141382 183454
rect 140826 182898 141062 183134
rect 141146 182898 141382 183134
rect 140826 147218 141062 147454
rect 141146 147218 141382 147454
rect 140826 146898 141062 147134
rect 141146 146898 141382 147134
rect 140826 111218 141062 111454
rect 141146 111218 141382 111454
rect 140826 110898 141062 111134
rect 141146 110898 141382 111134
rect 140826 75218 141062 75454
rect 141146 75218 141382 75454
rect 140826 74898 141062 75134
rect 141146 74898 141382 75134
rect 140826 39218 141062 39454
rect 141146 39218 141382 39454
rect 140826 38898 141062 39134
rect 141146 38898 141382 39134
rect 140826 3218 141062 3454
rect 141146 3218 141382 3454
rect 140826 2898 141062 3134
rect 141146 2898 141382 3134
rect 140826 -582 141062 -346
rect 141146 -582 141382 -346
rect 140826 -902 141062 -666
rect 141146 -902 141382 -666
rect 151986 710362 152222 710598
rect 152306 710362 152542 710598
rect 151986 710042 152222 710278
rect 152306 710042 152542 710278
rect 148266 708442 148502 708678
rect 148586 708442 148822 708678
rect 148266 708122 148502 708358
rect 148586 708122 148822 708358
rect 141986 680378 142222 680614
rect 142306 680378 142542 680614
rect 141986 680058 142222 680294
rect 142306 680058 142542 680294
rect 141986 644378 142222 644614
rect 142306 644378 142542 644614
rect 141986 644058 142222 644294
rect 142306 644058 142542 644294
rect 141986 608378 142222 608614
rect 142306 608378 142542 608614
rect 141986 608058 142222 608294
rect 142306 608058 142542 608294
rect 141986 572378 142222 572614
rect 142306 572378 142542 572614
rect 141986 572058 142222 572294
rect 142306 572058 142542 572294
rect 141986 536378 142222 536614
rect 142306 536378 142542 536614
rect 141986 536058 142222 536294
rect 142306 536058 142542 536294
rect 141986 500378 142222 500614
rect 142306 500378 142542 500614
rect 141986 500058 142222 500294
rect 142306 500058 142542 500294
rect 141986 464378 142222 464614
rect 142306 464378 142542 464614
rect 141986 464058 142222 464294
rect 142306 464058 142542 464294
rect 141986 428378 142222 428614
rect 142306 428378 142542 428614
rect 141986 428058 142222 428294
rect 142306 428058 142542 428294
rect 141986 392378 142222 392614
rect 142306 392378 142542 392614
rect 141986 392058 142222 392294
rect 142306 392058 142542 392294
rect 141986 356378 142222 356614
rect 142306 356378 142542 356614
rect 141986 356058 142222 356294
rect 142306 356058 142542 356294
rect 141986 320378 142222 320614
rect 142306 320378 142542 320614
rect 141986 320058 142222 320294
rect 142306 320058 142542 320294
rect 141986 284378 142222 284614
rect 142306 284378 142542 284614
rect 141986 284058 142222 284294
rect 142306 284058 142542 284294
rect 141986 248378 142222 248614
rect 142306 248378 142542 248614
rect 141986 248058 142222 248294
rect 142306 248058 142542 248294
rect 141986 212378 142222 212614
rect 142306 212378 142542 212614
rect 141986 212058 142222 212294
rect 142306 212058 142542 212294
rect 141986 176378 142222 176614
rect 142306 176378 142542 176614
rect 141986 176058 142222 176294
rect 142306 176058 142542 176294
rect 141986 140378 142222 140614
rect 142306 140378 142542 140614
rect 141986 140058 142222 140294
rect 142306 140058 142542 140294
rect 141986 104378 142222 104614
rect 142306 104378 142542 104614
rect 141986 104058 142222 104294
rect 142306 104058 142542 104294
rect 141986 68378 142222 68614
rect 142306 68378 142542 68614
rect 141986 68058 142222 68294
rect 142306 68058 142542 68294
rect 141986 32378 142222 32614
rect 142306 32378 142542 32614
rect 141986 32058 142222 32294
rect 142306 32058 142542 32294
rect 138266 -5382 138502 -5146
rect 138586 -5382 138822 -5146
rect 138266 -5702 138502 -5466
rect 138586 -5702 138822 -5466
rect 131986 -6342 132222 -6106
rect 132306 -6342 132542 -6106
rect 131986 -6662 132222 -6426
rect 132306 -6662 132542 -6426
rect 144546 706522 144782 706758
rect 144866 706522 145102 706758
rect 144546 706202 144782 706438
rect 144866 706202 145102 706438
rect 144546 690938 144782 691174
rect 144866 690938 145102 691174
rect 144546 690618 144782 690854
rect 144866 690618 145102 690854
rect 144546 654938 144782 655174
rect 144866 654938 145102 655174
rect 144546 654618 144782 654854
rect 144866 654618 145102 654854
rect 144546 618938 144782 619174
rect 144866 618938 145102 619174
rect 144546 618618 144782 618854
rect 144866 618618 145102 618854
rect 144546 582938 144782 583174
rect 144866 582938 145102 583174
rect 144546 582618 144782 582854
rect 144866 582618 145102 582854
rect 144546 546938 144782 547174
rect 144866 546938 145102 547174
rect 144546 546618 144782 546854
rect 144866 546618 145102 546854
rect 144546 510938 144782 511174
rect 144866 510938 145102 511174
rect 144546 510618 144782 510854
rect 144866 510618 145102 510854
rect 144546 474938 144782 475174
rect 144866 474938 145102 475174
rect 144546 474618 144782 474854
rect 144866 474618 145102 474854
rect 144546 438938 144782 439174
rect 144866 438938 145102 439174
rect 144546 438618 144782 438854
rect 144866 438618 145102 438854
rect 144546 402938 144782 403174
rect 144866 402938 145102 403174
rect 144546 402618 144782 402854
rect 144866 402618 145102 402854
rect 144546 366938 144782 367174
rect 144866 366938 145102 367174
rect 144546 366618 144782 366854
rect 144866 366618 145102 366854
rect 144546 330938 144782 331174
rect 144866 330938 145102 331174
rect 144546 330618 144782 330854
rect 144866 330618 145102 330854
rect 144546 294938 144782 295174
rect 144866 294938 145102 295174
rect 144546 294618 144782 294854
rect 144866 294618 145102 294854
rect 144546 258938 144782 259174
rect 144866 258938 145102 259174
rect 144546 258618 144782 258854
rect 144866 258618 145102 258854
rect 144546 222938 144782 223174
rect 144866 222938 145102 223174
rect 144546 222618 144782 222854
rect 144866 222618 145102 222854
rect 144546 186938 144782 187174
rect 144866 186938 145102 187174
rect 144546 186618 144782 186854
rect 144866 186618 145102 186854
rect 144546 150938 144782 151174
rect 144866 150938 145102 151174
rect 144546 150618 144782 150854
rect 144866 150618 145102 150854
rect 144546 114938 144782 115174
rect 144866 114938 145102 115174
rect 144546 114618 144782 114854
rect 144866 114618 145102 114854
rect 144546 78938 144782 79174
rect 144866 78938 145102 79174
rect 144546 78618 144782 78854
rect 144866 78618 145102 78854
rect 144546 42938 144782 43174
rect 144866 42938 145102 43174
rect 144546 42618 144782 42854
rect 144866 42618 145102 42854
rect 144546 6938 144782 7174
rect 144866 6938 145102 7174
rect 144546 6618 144782 6854
rect 144866 6618 145102 6854
rect 144546 -2502 144782 -2266
rect 144866 -2502 145102 -2266
rect 144546 -2822 144782 -2586
rect 144866 -2822 145102 -2586
rect 148266 694658 148502 694894
rect 148586 694658 148822 694894
rect 148266 694338 148502 694574
rect 148586 694338 148822 694574
rect 148266 658658 148502 658894
rect 148586 658658 148822 658894
rect 148266 658338 148502 658574
rect 148586 658338 148822 658574
rect 148266 622658 148502 622894
rect 148586 622658 148822 622894
rect 148266 622338 148502 622574
rect 148586 622338 148822 622574
rect 148266 586658 148502 586894
rect 148586 586658 148822 586894
rect 148266 586338 148502 586574
rect 148586 586338 148822 586574
rect 148266 550658 148502 550894
rect 148586 550658 148822 550894
rect 148266 550338 148502 550574
rect 148586 550338 148822 550574
rect 148266 514658 148502 514894
rect 148586 514658 148822 514894
rect 148266 514338 148502 514574
rect 148586 514338 148822 514574
rect 148266 478658 148502 478894
rect 148586 478658 148822 478894
rect 148266 478338 148502 478574
rect 148586 478338 148822 478574
rect 148266 442658 148502 442894
rect 148586 442658 148822 442894
rect 148266 442338 148502 442574
rect 148586 442338 148822 442574
rect 148266 406658 148502 406894
rect 148586 406658 148822 406894
rect 148266 406338 148502 406574
rect 148586 406338 148822 406574
rect 148266 370658 148502 370894
rect 148586 370658 148822 370894
rect 148266 370338 148502 370574
rect 148586 370338 148822 370574
rect 148266 334658 148502 334894
rect 148586 334658 148822 334894
rect 148266 334338 148502 334574
rect 148586 334338 148822 334574
rect 148266 298658 148502 298894
rect 148586 298658 148822 298894
rect 148266 298338 148502 298574
rect 148586 298338 148822 298574
rect 148266 262658 148502 262894
rect 148586 262658 148822 262894
rect 148266 262338 148502 262574
rect 148586 262338 148822 262574
rect 148266 226658 148502 226894
rect 148586 226658 148822 226894
rect 148266 226338 148502 226574
rect 148586 226338 148822 226574
rect 148266 190658 148502 190894
rect 148586 190658 148822 190894
rect 148266 190338 148502 190574
rect 148586 190338 148822 190574
rect 148266 154658 148502 154894
rect 148586 154658 148822 154894
rect 148266 154338 148502 154574
rect 148586 154338 148822 154574
rect 148266 118658 148502 118894
rect 148586 118658 148822 118894
rect 148266 118338 148502 118574
rect 148586 118338 148822 118574
rect 148266 82658 148502 82894
rect 148586 82658 148822 82894
rect 148266 82338 148502 82574
rect 148586 82338 148822 82574
rect 148266 46658 148502 46894
rect 148586 46658 148822 46894
rect 148266 46338 148502 46574
rect 148586 46338 148822 46574
rect 148266 10658 148502 10894
rect 148586 10658 148822 10894
rect 148266 10338 148502 10574
rect 148586 10338 148822 10574
rect 150826 705562 151062 705798
rect 151146 705562 151382 705798
rect 150826 705242 151062 705478
rect 151146 705242 151382 705478
rect 150826 669218 151062 669454
rect 151146 669218 151382 669454
rect 150826 668898 151062 669134
rect 151146 668898 151382 669134
rect 150826 633218 151062 633454
rect 151146 633218 151382 633454
rect 150826 632898 151062 633134
rect 151146 632898 151382 633134
rect 150826 597218 151062 597454
rect 151146 597218 151382 597454
rect 150826 596898 151062 597134
rect 151146 596898 151382 597134
rect 150826 561218 151062 561454
rect 151146 561218 151382 561454
rect 150826 560898 151062 561134
rect 151146 560898 151382 561134
rect 150826 525218 151062 525454
rect 151146 525218 151382 525454
rect 150826 524898 151062 525134
rect 151146 524898 151382 525134
rect 150826 489218 151062 489454
rect 151146 489218 151382 489454
rect 150826 488898 151062 489134
rect 151146 488898 151382 489134
rect 150826 453218 151062 453454
rect 151146 453218 151382 453454
rect 150826 452898 151062 453134
rect 151146 452898 151382 453134
rect 150826 417218 151062 417454
rect 151146 417218 151382 417454
rect 150826 416898 151062 417134
rect 151146 416898 151382 417134
rect 150826 381218 151062 381454
rect 151146 381218 151382 381454
rect 150826 380898 151062 381134
rect 151146 380898 151382 381134
rect 150826 345218 151062 345454
rect 151146 345218 151382 345454
rect 150826 344898 151062 345134
rect 151146 344898 151382 345134
rect 150826 309218 151062 309454
rect 151146 309218 151382 309454
rect 150826 308898 151062 309134
rect 151146 308898 151382 309134
rect 150826 273218 151062 273454
rect 151146 273218 151382 273454
rect 150826 272898 151062 273134
rect 151146 272898 151382 273134
rect 150826 237218 151062 237454
rect 151146 237218 151382 237454
rect 150826 236898 151062 237134
rect 151146 236898 151382 237134
rect 150826 201218 151062 201454
rect 151146 201218 151382 201454
rect 150826 200898 151062 201134
rect 151146 200898 151382 201134
rect 150826 165218 151062 165454
rect 151146 165218 151382 165454
rect 150826 164898 151062 165134
rect 151146 164898 151382 165134
rect 150826 129218 151062 129454
rect 151146 129218 151382 129454
rect 150826 128898 151062 129134
rect 151146 128898 151382 129134
rect 150826 93218 151062 93454
rect 151146 93218 151382 93454
rect 150826 92898 151062 93134
rect 151146 92898 151382 93134
rect 150826 57218 151062 57454
rect 151146 57218 151382 57454
rect 150826 56898 151062 57134
rect 151146 56898 151382 57134
rect 150826 21218 151062 21454
rect 151146 21218 151382 21454
rect 150826 20898 151062 21134
rect 151146 20898 151382 21134
rect 150826 -1542 151062 -1306
rect 151146 -1542 151382 -1306
rect 150826 -1862 151062 -1626
rect 151146 -1862 151382 -1626
rect 161986 711322 162222 711558
rect 162306 711322 162542 711558
rect 161986 711002 162222 711238
rect 162306 711002 162542 711238
rect 158266 709402 158502 709638
rect 158586 709402 158822 709638
rect 158266 709082 158502 709318
rect 158586 709082 158822 709318
rect 151986 698378 152222 698614
rect 152306 698378 152542 698614
rect 151986 698058 152222 698294
rect 152306 698058 152542 698294
rect 151986 662378 152222 662614
rect 152306 662378 152542 662614
rect 151986 662058 152222 662294
rect 152306 662058 152542 662294
rect 151986 626378 152222 626614
rect 152306 626378 152542 626614
rect 151986 626058 152222 626294
rect 152306 626058 152542 626294
rect 151986 590378 152222 590614
rect 152306 590378 152542 590614
rect 151986 590058 152222 590294
rect 152306 590058 152542 590294
rect 151986 554378 152222 554614
rect 152306 554378 152542 554614
rect 151986 554058 152222 554294
rect 152306 554058 152542 554294
rect 151986 518378 152222 518614
rect 152306 518378 152542 518614
rect 151986 518058 152222 518294
rect 152306 518058 152542 518294
rect 151986 482378 152222 482614
rect 152306 482378 152542 482614
rect 151986 482058 152222 482294
rect 152306 482058 152542 482294
rect 151986 446378 152222 446614
rect 152306 446378 152542 446614
rect 151986 446058 152222 446294
rect 152306 446058 152542 446294
rect 151986 410378 152222 410614
rect 152306 410378 152542 410614
rect 151986 410058 152222 410294
rect 152306 410058 152542 410294
rect 151986 374378 152222 374614
rect 152306 374378 152542 374614
rect 151986 374058 152222 374294
rect 152306 374058 152542 374294
rect 151986 338378 152222 338614
rect 152306 338378 152542 338614
rect 151986 338058 152222 338294
rect 152306 338058 152542 338294
rect 151986 302378 152222 302614
rect 152306 302378 152542 302614
rect 151986 302058 152222 302294
rect 152306 302058 152542 302294
rect 151986 266378 152222 266614
rect 152306 266378 152542 266614
rect 151986 266058 152222 266294
rect 152306 266058 152542 266294
rect 151986 230378 152222 230614
rect 152306 230378 152542 230614
rect 151986 230058 152222 230294
rect 152306 230058 152542 230294
rect 151986 194378 152222 194614
rect 152306 194378 152542 194614
rect 151986 194058 152222 194294
rect 152306 194058 152542 194294
rect 151986 158378 152222 158614
rect 152306 158378 152542 158614
rect 151986 158058 152222 158294
rect 152306 158058 152542 158294
rect 151986 122378 152222 122614
rect 152306 122378 152542 122614
rect 151986 122058 152222 122294
rect 152306 122058 152542 122294
rect 151986 86378 152222 86614
rect 152306 86378 152542 86614
rect 151986 86058 152222 86294
rect 152306 86058 152542 86294
rect 151986 50378 152222 50614
rect 152306 50378 152542 50614
rect 151986 50058 152222 50294
rect 152306 50058 152542 50294
rect 151986 14378 152222 14614
rect 152306 14378 152542 14614
rect 151986 14058 152222 14294
rect 152306 14058 152542 14294
rect 148266 -4422 148502 -4186
rect 148586 -4422 148822 -4186
rect 148266 -4742 148502 -4506
rect 148586 -4742 148822 -4506
rect 141986 -7302 142222 -7066
rect 142306 -7302 142542 -7066
rect 141986 -7622 142222 -7386
rect 142306 -7622 142542 -7386
rect 154546 707482 154782 707718
rect 154866 707482 155102 707718
rect 154546 707162 154782 707398
rect 154866 707162 155102 707398
rect 154546 672938 154782 673174
rect 154866 672938 155102 673174
rect 154546 672618 154782 672854
rect 154866 672618 155102 672854
rect 154546 636938 154782 637174
rect 154866 636938 155102 637174
rect 154546 636618 154782 636854
rect 154866 636618 155102 636854
rect 154546 600938 154782 601174
rect 154866 600938 155102 601174
rect 154546 600618 154782 600854
rect 154866 600618 155102 600854
rect 154546 564938 154782 565174
rect 154866 564938 155102 565174
rect 154546 564618 154782 564854
rect 154866 564618 155102 564854
rect 154546 528938 154782 529174
rect 154866 528938 155102 529174
rect 154546 528618 154782 528854
rect 154866 528618 155102 528854
rect 154546 492938 154782 493174
rect 154866 492938 155102 493174
rect 154546 492618 154782 492854
rect 154866 492618 155102 492854
rect 154546 456938 154782 457174
rect 154866 456938 155102 457174
rect 154546 456618 154782 456854
rect 154866 456618 155102 456854
rect 154546 420938 154782 421174
rect 154866 420938 155102 421174
rect 154546 420618 154782 420854
rect 154866 420618 155102 420854
rect 154546 384938 154782 385174
rect 154866 384938 155102 385174
rect 154546 384618 154782 384854
rect 154866 384618 155102 384854
rect 154546 348938 154782 349174
rect 154866 348938 155102 349174
rect 154546 348618 154782 348854
rect 154866 348618 155102 348854
rect 154546 312938 154782 313174
rect 154866 312938 155102 313174
rect 154546 312618 154782 312854
rect 154866 312618 155102 312854
rect 154546 276938 154782 277174
rect 154866 276938 155102 277174
rect 154546 276618 154782 276854
rect 154866 276618 155102 276854
rect 154546 240938 154782 241174
rect 154866 240938 155102 241174
rect 154546 240618 154782 240854
rect 154866 240618 155102 240854
rect 154546 204938 154782 205174
rect 154866 204938 155102 205174
rect 154546 204618 154782 204854
rect 154866 204618 155102 204854
rect 154546 168938 154782 169174
rect 154866 168938 155102 169174
rect 154546 168618 154782 168854
rect 154866 168618 155102 168854
rect 154546 132938 154782 133174
rect 154866 132938 155102 133174
rect 154546 132618 154782 132854
rect 154866 132618 155102 132854
rect 154546 96938 154782 97174
rect 154866 96938 155102 97174
rect 154546 96618 154782 96854
rect 154866 96618 155102 96854
rect 154546 60938 154782 61174
rect 154866 60938 155102 61174
rect 154546 60618 154782 60854
rect 154866 60618 155102 60854
rect 154546 24938 154782 25174
rect 154866 24938 155102 25174
rect 154546 24618 154782 24854
rect 154866 24618 155102 24854
rect 154546 -3462 154782 -3226
rect 154866 -3462 155102 -3226
rect 154546 -3782 154782 -3546
rect 154866 -3782 155102 -3546
rect 158266 676658 158502 676894
rect 158586 676658 158822 676894
rect 158266 676338 158502 676574
rect 158586 676338 158822 676574
rect 158266 640658 158502 640894
rect 158586 640658 158822 640894
rect 158266 640338 158502 640574
rect 158586 640338 158822 640574
rect 158266 604658 158502 604894
rect 158586 604658 158822 604894
rect 158266 604338 158502 604574
rect 158586 604338 158822 604574
rect 158266 568658 158502 568894
rect 158586 568658 158822 568894
rect 158266 568338 158502 568574
rect 158586 568338 158822 568574
rect 158266 532658 158502 532894
rect 158586 532658 158822 532894
rect 158266 532338 158502 532574
rect 158586 532338 158822 532574
rect 158266 496658 158502 496894
rect 158586 496658 158822 496894
rect 158266 496338 158502 496574
rect 158586 496338 158822 496574
rect 158266 460658 158502 460894
rect 158586 460658 158822 460894
rect 158266 460338 158502 460574
rect 158586 460338 158822 460574
rect 158266 424658 158502 424894
rect 158586 424658 158822 424894
rect 158266 424338 158502 424574
rect 158586 424338 158822 424574
rect 158266 388658 158502 388894
rect 158586 388658 158822 388894
rect 158266 388338 158502 388574
rect 158586 388338 158822 388574
rect 158266 352658 158502 352894
rect 158586 352658 158822 352894
rect 158266 352338 158502 352574
rect 158586 352338 158822 352574
rect 158266 316658 158502 316894
rect 158586 316658 158822 316894
rect 158266 316338 158502 316574
rect 158586 316338 158822 316574
rect 158266 280658 158502 280894
rect 158586 280658 158822 280894
rect 158266 280338 158502 280574
rect 158586 280338 158822 280574
rect 158266 244658 158502 244894
rect 158586 244658 158822 244894
rect 158266 244338 158502 244574
rect 158586 244338 158822 244574
rect 158266 208658 158502 208894
rect 158586 208658 158822 208894
rect 158266 208338 158502 208574
rect 158586 208338 158822 208574
rect 158266 172658 158502 172894
rect 158586 172658 158822 172894
rect 158266 172338 158502 172574
rect 158586 172338 158822 172574
rect 158266 136658 158502 136894
rect 158586 136658 158822 136894
rect 158266 136338 158502 136574
rect 158586 136338 158822 136574
rect 158266 100658 158502 100894
rect 158586 100658 158822 100894
rect 158266 100338 158502 100574
rect 158586 100338 158822 100574
rect 158266 64658 158502 64894
rect 158586 64658 158822 64894
rect 158266 64338 158502 64574
rect 158586 64338 158822 64574
rect 158266 28658 158502 28894
rect 158586 28658 158822 28894
rect 158266 28338 158502 28574
rect 158586 28338 158822 28574
rect 160826 704602 161062 704838
rect 161146 704602 161382 704838
rect 160826 704282 161062 704518
rect 161146 704282 161382 704518
rect 160826 687218 161062 687454
rect 161146 687218 161382 687454
rect 160826 686898 161062 687134
rect 161146 686898 161382 687134
rect 160826 651218 161062 651454
rect 161146 651218 161382 651454
rect 160826 650898 161062 651134
rect 161146 650898 161382 651134
rect 160826 615218 161062 615454
rect 161146 615218 161382 615454
rect 160826 614898 161062 615134
rect 161146 614898 161382 615134
rect 160826 579218 161062 579454
rect 161146 579218 161382 579454
rect 160826 578898 161062 579134
rect 161146 578898 161382 579134
rect 160826 543218 161062 543454
rect 161146 543218 161382 543454
rect 160826 542898 161062 543134
rect 161146 542898 161382 543134
rect 160826 507218 161062 507454
rect 161146 507218 161382 507454
rect 160826 506898 161062 507134
rect 161146 506898 161382 507134
rect 160826 471218 161062 471454
rect 161146 471218 161382 471454
rect 160826 470898 161062 471134
rect 161146 470898 161382 471134
rect 160826 435218 161062 435454
rect 161146 435218 161382 435454
rect 160826 434898 161062 435134
rect 161146 434898 161382 435134
rect 160826 399218 161062 399454
rect 161146 399218 161382 399454
rect 160826 398898 161062 399134
rect 161146 398898 161382 399134
rect 160826 363218 161062 363454
rect 161146 363218 161382 363454
rect 160826 362898 161062 363134
rect 161146 362898 161382 363134
rect 160826 327218 161062 327454
rect 161146 327218 161382 327454
rect 160826 326898 161062 327134
rect 161146 326898 161382 327134
rect 160826 291218 161062 291454
rect 161146 291218 161382 291454
rect 160826 290898 161062 291134
rect 161146 290898 161382 291134
rect 160826 255218 161062 255454
rect 161146 255218 161382 255454
rect 160826 254898 161062 255134
rect 161146 254898 161382 255134
rect 160826 219218 161062 219454
rect 161146 219218 161382 219454
rect 160826 218898 161062 219134
rect 161146 218898 161382 219134
rect 160826 183218 161062 183454
rect 161146 183218 161382 183454
rect 160826 182898 161062 183134
rect 161146 182898 161382 183134
rect 160826 147218 161062 147454
rect 161146 147218 161382 147454
rect 160826 146898 161062 147134
rect 161146 146898 161382 147134
rect 160826 111218 161062 111454
rect 161146 111218 161382 111454
rect 160826 110898 161062 111134
rect 161146 110898 161382 111134
rect 160826 75218 161062 75454
rect 161146 75218 161382 75454
rect 160826 74898 161062 75134
rect 161146 74898 161382 75134
rect 160826 39218 161062 39454
rect 161146 39218 161382 39454
rect 160826 38898 161062 39134
rect 161146 38898 161382 39134
rect 160826 3218 161062 3454
rect 161146 3218 161382 3454
rect 160826 2898 161062 3134
rect 161146 2898 161382 3134
rect 160826 -582 161062 -346
rect 161146 -582 161382 -346
rect 160826 -902 161062 -666
rect 161146 -902 161382 -666
rect 171986 710362 172222 710598
rect 172306 710362 172542 710598
rect 171986 710042 172222 710278
rect 172306 710042 172542 710278
rect 168266 708442 168502 708678
rect 168586 708442 168822 708678
rect 168266 708122 168502 708358
rect 168586 708122 168822 708358
rect 161986 680378 162222 680614
rect 162306 680378 162542 680614
rect 161986 680058 162222 680294
rect 162306 680058 162542 680294
rect 161986 644378 162222 644614
rect 162306 644378 162542 644614
rect 161986 644058 162222 644294
rect 162306 644058 162542 644294
rect 161986 608378 162222 608614
rect 162306 608378 162542 608614
rect 161986 608058 162222 608294
rect 162306 608058 162542 608294
rect 161986 572378 162222 572614
rect 162306 572378 162542 572614
rect 161986 572058 162222 572294
rect 162306 572058 162542 572294
rect 161986 536378 162222 536614
rect 162306 536378 162542 536614
rect 161986 536058 162222 536294
rect 162306 536058 162542 536294
rect 161986 500378 162222 500614
rect 162306 500378 162542 500614
rect 161986 500058 162222 500294
rect 162306 500058 162542 500294
rect 161986 464378 162222 464614
rect 162306 464378 162542 464614
rect 161986 464058 162222 464294
rect 162306 464058 162542 464294
rect 161986 428378 162222 428614
rect 162306 428378 162542 428614
rect 161986 428058 162222 428294
rect 162306 428058 162542 428294
rect 161986 392378 162222 392614
rect 162306 392378 162542 392614
rect 161986 392058 162222 392294
rect 162306 392058 162542 392294
rect 161986 356378 162222 356614
rect 162306 356378 162542 356614
rect 161986 356058 162222 356294
rect 162306 356058 162542 356294
rect 161986 320378 162222 320614
rect 162306 320378 162542 320614
rect 161986 320058 162222 320294
rect 162306 320058 162542 320294
rect 161986 284378 162222 284614
rect 162306 284378 162542 284614
rect 161986 284058 162222 284294
rect 162306 284058 162542 284294
rect 161986 248378 162222 248614
rect 162306 248378 162542 248614
rect 161986 248058 162222 248294
rect 162306 248058 162542 248294
rect 161986 212378 162222 212614
rect 162306 212378 162542 212614
rect 161986 212058 162222 212294
rect 162306 212058 162542 212294
rect 161986 176378 162222 176614
rect 162306 176378 162542 176614
rect 161986 176058 162222 176294
rect 162306 176058 162542 176294
rect 161986 140378 162222 140614
rect 162306 140378 162542 140614
rect 161986 140058 162222 140294
rect 162306 140058 162542 140294
rect 161986 104378 162222 104614
rect 162306 104378 162542 104614
rect 161986 104058 162222 104294
rect 162306 104058 162542 104294
rect 161986 68378 162222 68614
rect 162306 68378 162542 68614
rect 161986 68058 162222 68294
rect 162306 68058 162542 68294
rect 161986 32378 162222 32614
rect 162306 32378 162542 32614
rect 161986 32058 162222 32294
rect 162306 32058 162542 32294
rect 158266 -5382 158502 -5146
rect 158586 -5382 158822 -5146
rect 158266 -5702 158502 -5466
rect 158586 -5702 158822 -5466
rect 151986 -6342 152222 -6106
rect 152306 -6342 152542 -6106
rect 151986 -6662 152222 -6426
rect 152306 -6662 152542 -6426
rect 164546 706522 164782 706758
rect 164866 706522 165102 706758
rect 164546 706202 164782 706438
rect 164866 706202 165102 706438
rect 164546 690938 164782 691174
rect 164866 690938 165102 691174
rect 164546 690618 164782 690854
rect 164866 690618 165102 690854
rect 164546 654938 164782 655174
rect 164866 654938 165102 655174
rect 164546 654618 164782 654854
rect 164866 654618 165102 654854
rect 164546 618938 164782 619174
rect 164866 618938 165102 619174
rect 164546 618618 164782 618854
rect 164866 618618 165102 618854
rect 164546 582938 164782 583174
rect 164866 582938 165102 583174
rect 164546 582618 164782 582854
rect 164866 582618 165102 582854
rect 164546 546938 164782 547174
rect 164866 546938 165102 547174
rect 164546 546618 164782 546854
rect 164866 546618 165102 546854
rect 164546 510938 164782 511174
rect 164866 510938 165102 511174
rect 164546 510618 164782 510854
rect 164866 510618 165102 510854
rect 164546 474938 164782 475174
rect 164866 474938 165102 475174
rect 164546 474618 164782 474854
rect 164866 474618 165102 474854
rect 164546 438938 164782 439174
rect 164866 438938 165102 439174
rect 164546 438618 164782 438854
rect 164866 438618 165102 438854
rect 164546 402938 164782 403174
rect 164866 402938 165102 403174
rect 164546 402618 164782 402854
rect 164866 402618 165102 402854
rect 164546 366938 164782 367174
rect 164866 366938 165102 367174
rect 164546 366618 164782 366854
rect 164866 366618 165102 366854
rect 164546 330938 164782 331174
rect 164866 330938 165102 331174
rect 164546 330618 164782 330854
rect 164866 330618 165102 330854
rect 164546 294938 164782 295174
rect 164866 294938 165102 295174
rect 164546 294618 164782 294854
rect 164866 294618 165102 294854
rect 164546 258938 164782 259174
rect 164866 258938 165102 259174
rect 164546 258618 164782 258854
rect 164866 258618 165102 258854
rect 164546 222938 164782 223174
rect 164866 222938 165102 223174
rect 164546 222618 164782 222854
rect 164866 222618 165102 222854
rect 164546 186938 164782 187174
rect 164866 186938 165102 187174
rect 164546 186618 164782 186854
rect 164866 186618 165102 186854
rect 164546 150938 164782 151174
rect 164866 150938 165102 151174
rect 164546 150618 164782 150854
rect 164866 150618 165102 150854
rect 164546 114938 164782 115174
rect 164866 114938 165102 115174
rect 164546 114618 164782 114854
rect 164866 114618 165102 114854
rect 164546 78938 164782 79174
rect 164866 78938 165102 79174
rect 164546 78618 164782 78854
rect 164866 78618 165102 78854
rect 164546 42938 164782 43174
rect 164866 42938 165102 43174
rect 164546 42618 164782 42854
rect 164866 42618 165102 42854
rect 164546 6938 164782 7174
rect 164866 6938 165102 7174
rect 164546 6618 164782 6854
rect 164866 6618 165102 6854
rect 164546 -2502 164782 -2266
rect 164866 -2502 165102 -2266
rect 164546 -2822 164782 -2586
rect 164866 -2822 165102 -2586
rect 168266 694658 168502 694894
rect 168586 694658 168822 694894
rect 168266 694338 168502 694574
rect 168586 694338 168822 694574
rect 168266 658658 168502 658894
rect 168586 658658 168822 658894
rect 168266 658338 168502 658574
rect 168586 658338 168822 658574
rect 168266 622658 168502 622894
rect 168586 622658 168822 622894
rect 168266 622338 168502 622574
rect 168586 622338 168822 622574
rect 168266 586658 168502 586894
rect 168586 586658 168822 586894
rect 168266 586338 168502 586574
rect 168586 586338 168822 586574
rect 168266 550658 168502 550894
rect 168586 550658 168822 550894
rect 168266 550338 168502 550574
rect 168586 550338 168822 550574
rect 168266 514658 168502 514894
rect 168586 514658 168822 514894
rect 168266 514338 168502 514574
rect 168586 514338 168822 514574
rect 168266 478658 168502 478894
rect 168586 478658 168822 478894
rect 168266 478338 168502 478574
rect 168586 478338 168822 478574
rect 168266 442658 168502 442894
rect 168586 442658 168822 442894
rect 168266 442338 168502 442574
rect 168586 442338 168822 442574
rect 168266 406658 168502 406894
rect 168586 406658 168822 406894
rect 168266 406338 168502 406574
rect 168586 406338 168822 406574
rect 168266 370658 168502 370894
rect 168586 370658 168822 370894
rect 168266 370338 168502 370574
rect 168586 370338 168822 370574
rect 168266 334658 168502 334894
rect 168586 334658 168822 334894
rect 168266 334338 168502 334574
rect 168586 334338 168822 334574
rect 168266 298658 168502 298894
rect 168586 298658 168822 298894
rect 168266 298338 168502 298574
rect 168586 298338 168822 298574
rect 168266 262658 168502 262894
rect 168586 262658 168822 262894
rect 168266 262338 168502 262574
rect 168586 262338 168822 262574
rect 168266 226658 168502 226894
rect 168586 226658 168822 226894
rect 168266 226338 168502 226574
rect 168586 226338 168822 226574
rect 168266 190658 168502 190894
rect 168586 190658 168822 190894
rect 168266 190338 168502 190574
rect 168586 190338 168822 190574
rect 168266 154658 168502 154894
rect 168586 154658 168822 154894
rect 168266 154338 168502 154574
rect 168586 154338 168822 154574
rect 168266 118658 168502 118894
rect 168586 118658 168822 118894
rect 168266 118338 168502 118574
rect 168586 118338 168822 118574
rect 168266 82658 168502 82894
rect 168586 82658 168822 82894
rect 168266 82338 168502 82574
rect 168586 82338 168822 82574
rect 168266 46658 168502 46894
rect 168586 46658 168822 46894
rect 168266 46338 168502 46574
rect 168586 46338 168822 46574
rect 168266 10658 168502 10894
rect 168586 10658 168822 10894
rect 168266 10338 168502 10574
rect 168586 10338 168822 10574
rect 170826 705562 171062 705798
rect 171146 705562 171382 705798
rect 170826 705242 171062 705478
rect 171146 705242 171382 705478
rect 170826 669218 171062 669454
rect 171146 669218 171382 669454
rect 170826 668898 171062 669134
rect 171146 668898 171382 669134
rect 170826 633218 171062 633454
rect 171146 633218 171382 633454
rect 170826 632898 171062 633134
rect 171146 632898 171382 633134
rect 170826 597218 171062 597454
rect 171146 597218 171382 597454
rect 170826 596898 171062 597134
rect 171146 596898 171382 597134
rect 170826 561218 171062 561454
rect 171146 561218 171382 561454
rect 170826 560898 171062 561134
rect 171146 560898 171382 561134
rect 170826 525218 171062 525454
rect 171146 525218 171382 525454
rect 170826 524898 171062 525134
rect 171146 524898 171382 525134
rect 170826 489218 171062 489454
rect 171146 489218 171382 489454
rect 170826 488898 171062 489134
rect 171146 488898 171382 489134
rect 170826 453218 171062 453454
rect 171146 453218 171382 453454
rect 170826 452898 171062 453134
rect 171146 452898 171382 453134
rect 170826 417218 171062 417454
rect 171146 417218 171382 417454
rect 170826 416898 171062 417134
rect 171146 416898 171382 417134
rect 170826 381218 171062 381454
rect 171146 381218 171382 381454
rect 170826 380898 171062 381134
rect 171146 380898 171382 381134
rect 170826 345218 171062 345454
rect 171146 345218 171382 345454
rect 170826 344898 171062 345134
rect 171146 344898 171382 345134
rect 170826 309218 171062 309454
rect 171146 309218 171382 309454
rect 170826 308898 171062 309134
rect 171146 308898 171382 309134
rect 170826 273218 171062 273454
rect 171146 273218 171382 273454
rect 170826 272898 171062 273134
rect 171146 272898 171382 273134
rect 170826 237218 171062 237454
rect 171146 237218 171382 237454
rect 170826 236898 171062 237134
rect 171146 236898 171382 237134
rect 170826 201218 171062 201454
rect 171146 201218 171382 201454
rect 170826 200898 171062 201134
rect 171146 200898 171382 201134
rect 170826 165218 171062 165454
rect 171146 165218 171382 165454
rect 170826 164898 171062 165134
rect 171146 164898 171382 165134
rect 170826 129218 171062 129454
rect 171146 129218 171382 129454
rect 170826 128898 171062 129134
rect 171146 128898 171382 129134
rect 170826 93218 171062 93454
rect 171146 93218 171382 93454
rect 170826 92898 171062 93134
rect 171146 92898 171382 93134
rect 170826 57218 171062 57454
rect 171146 57218 171382 57454
rect 170826 56898 171062 57134
rect 171146 56898 171382 57134
rect 170826 21218 171062 21454
rect 171146 21218 171382 21454
rect 170826 20898 171062 21134
rect 171146 20898 171382 21134
rect 170826 -1542 171062 -1306
rect 171146 -1542 171382 -1306
rect 170826 -1862 171062 -1626
rect 171146 -1862 171382 -1626
rect 181986 711322 182222 711558
rect 182306 711322 182542 711558
rect 181986 711002 182222 711238
rect 182306 711002 182542 711238
rect 178266 709402 178502 709638
rect 178586 709402 178822 709638
rect 178266 709082 178502 709318
rect 178586 709082 178822 709318
rect 171986 698378 172222 698614
rect 172306 698378 172542 698614
rect 171986 698058 172222 698294
rect 172306 698058 172542 698294
rect 171986 662378 172222 662614
rect 172306 662378 172542 662614
rect 171986 662058 172222 662294
rect 172306 662058 172542 662294
rect 171986 626378 172222 626614
rect 172306 626378 172542 626614
rect 171986 626058 172222 626294
rect 172306 626058 172542 626294
rect 171986 590378 172222 590614
rect 172306 590378 172542 590614
rect 171986 590058 172222 590294
rect 172306 590058 172542 590294
rect 171986 554378 172222 554614
rect 172306 554378 172542 554614
rect 171986 554058 172222 554294
rect 172306 554058 172542 554294
rect 171986 518378 172222 518614
rect 172306 518378 172542 518614
rect 171986 518058 172222 518294
rect 172306 518058 172542 518294
rect 171986 482378 172222 482614
rect 172306 482378 172542 482614
rect 171986 482058 172222 482294
rect 172306 482058 172542 482294
rect 171986 446378 172222 446614
rect 172306 446378 172542 446614
rect 171986 446058 172222 446294
rect 172306 446058 172542 446294
rect 171986 410378 172222 410614
rect 172306 410378 172542 410614
rect 171986 410058 172222 410294
rect 172306 410058 172542 410294
rect 171986 374378 172222 374614
rect 172306 374378 172542 374614
rect 171986 374058 172222 374294
rect 172306 374058 172542 374294
rect 171986 338378 172222 338614
rect 172306 338378 172542 338614
rect 171986 338058 172222 338294
rect 172306 338058 172542 338294
rect 171986 302378 172222 302614
rect 172306 302378 172542 302614
rect 171986 302058 172222 302294
rect 172306 302058 172542 302294
rect 171986 266378 172222 266614
rect 172306 266378 172542 266614
rect 171986 266058 172222 266294
rect 172306 266058 172542 266294
rect 171986 230378 172222 230614
rect 172306 230378 172542 230614
rect 171986 230058 172222 230294
rect 172306 230058 172542 230294
rect 171986 194378 172222 194614
rect 172306 194378 172542 194614
rect 171986 194058 172222 194294
rect 172306 194058 172542 194294
rect 171986 158378 172222 158614
rect 172306 158378 172542 158614
rect 171986 158058 172222 158294
rect 172306 158058 172542 158294
rect 171986 122378 172222 122614
rect 172306 122378 172542 122614
rect 171986 122058 172222 122294
rect 172306 122058 172542 122294
rect 171986 86378 172222 86614
rect 172306 86378 172542 86614
rect 171986 86058 172222 86294
rect 172306 86058 172542 86294
rect 171986 50378 172222 50614
rect 172306 50378 172542 50614
rect 171986 50058 172222 50294
rect 172306 50058 172542 50294
rect 171986 14378 172222 14614
rect 172306 14378 172542 14614
rect 171986 14058 172222 14294
rect 172306 14058 172542 14294
rect 168266 -4422 168502 -4186
rect 168586 -4422 168822 -4186
rect 168266 -4742 168502 -4506
rect 168586 -4742 168822 -4506
rect 161986 -7302 162222 -7066
rect 162306 -7302 162542 -7066
rect 161986 -7622 162222 -7386
rect 162306 -7622 162542 -7386
rect 174546 707482 174782 707718
rect 174866 707482 175102 707718
rect 174546 707162 174782 707398
rect 174866 707162 175102 707398
rect 174546 672938 174782 673174
rect 174866 672938 175102 673174
rect 174546 672618 174782 672854
rect 174866 672618 175102 672854
rect 174546 636938 174782 637174
rect 174866 636938 175102 637174
rect 174546 636618 174782 636854
rect 174866 636618 175102 636854
rect 174546 600938 174782 601174
rect 174866 600938 175102 601174
rect 174546 600618 174782 600854
rect 174866 600618 175102 600854
rect 174546 564938 174782 565174
rect 174866 564938 175102 565174
rect 174546 564618 174782 564854
rect 174866 564618 175102 564854
rect 174546 528938 174782 529174
rect 174866 528938 175102 529174
rect 174546 528618 174782 528854
rect 174866 528618 175102 528854
rect 174546 492938 174782 493174
rect 174866 492938 175102 493174
rect 174546 492618 174782 492854
rect 174866 492618 175102 492854
rect 174546 456938 174782 457174
rect 174866 456938 175102 457174
rect 174546 456618 174782 456854
rect 174866 456618 175102 456854
rect 174546 420938 174782 421174
rect 174866 420938 175102 421174
rect 174546 420618 174782 420854
rect 174866 420618 175102 420854
rect 174546 384938 174782 385174
rect 174866 384938 175102 385174
rect 174546 384618 174782 384854
rect 174866 384618 175102 384854
rect 174546 348938 174782 349174
rect 174866 348938 175102 349174
rect 174546 348618 174782 348854
rect 174866 348618 175102 348854
rect 174546 312938 174782 313174
rect 174866 312938 175102 313174
rect 174546 312618 174782 312854
rect 174866 312618 175102 312854
rect 174546 276938 174782 277174
rect 174866 276938 175102 277174
rect 174546 276618 174782 276854
rect 174866 276618 175102 276854
rect 174546 240938 174782 241174
rect 174866 240938 175102 241174
rect 174546 240618 174782 240854
rect 174866 240618 175102 240854
rect 174546 204938 174782 205174
rect 174866 204938 175102 205174
rect 174546 204618 174782 204854
rect 174866 204618 175102 204854
rect 174546 168938 174782 169174
rect 174866 168938 175102 169174
rect 174546 168618 174782 168854
rect 174866 168618 175102 168854
rect 174546 132938 174782 133174
rect 174866 132938 175102 133174
rect 174546 132618 174782 132854
rect 174866 132618 175102 132854
rect 174546 96938 174782 97174
rect 174866 96938 175102 97174
rect 174546 96618 174782 96854
rect 174866 96618 175102 96854
rect 174546 60938 174782 61174
rect 174866 60938 175102 61174
rect 174546 60618 174782 60854
rect 174866 60618 175102 60854
rect 174546 24938 174782 25174
rect 174866 24938 175102 25174
rect 174546 24618 174782 24854
rect 174866 24618 175102 24854
rect 174546 -3462 174782 -3226
rect 174866 -3462 175102 -3226
rect 174546 -3782 174782 -3546
rect 174866 -3782 175102 -3546
rect 178266 676658 178502 676894
rect 178586 676658 178822 676894
rect 178266 676338 178502 676574
rect 178586 676338 178822 676574
rect 178266 640658 178502 640894
rect 178586 640658 178822 640894
rect 178266 640338 178502 640574
rect 178586 640338 178822 640574
rect 178266 604658 178502 604894
rect 178586 604658 178822 604894
rect 178266 604338 178502 604574
rect 178586 604338 178822 604574
rect 178266 568658 178502 568894
rect 178586 568658 178822 568894
rect 178266 568338 178502 568574
rect 178586 568338 178822 568574
rect 178266 532658 178502 532894
rect 178586 532658 178822 532894
rect 178266 532338 178502 532574
rect 178586 532338 178822 532574
rect 178266 496658 178502 496894
rect 178586 496658 178822 496894
rect 178266 496338 178502 496574
rect 178586 496338 178822 496574
rect 178266 460658 178502 460894
rect 178586 460658 178822 460894
rect 178266 460338 178502 460574
rect 178586 460338 178822 460574
rect 178266 424658 178502 424894
rect 178586 424658 178822 424894
rect 178266 424338 178502 424574
rect 178586 424338 178822 424574
rect 178266 388658 178502 388894
rect 178586 388658 178822 388894
rect 178266 388338 178502 388574
rect 178586 388338 178822 388574
rect 178266 352658 178502 352894
rect 178586 352658 178822 352894
rect 178266 352338 178502 352574
rect 178586 352338 178822 352574
rect 178266 316658 178502 316894
rect 178586 316658 178822 316894
rect 178266 316338 178502 316574
rect 178586 316338 178822 316574
rect 178266 280658 178502 280894
rect 178586 280658 178822 280894
rect 178266 280338 178502 280574
rect 178586 280338 178822 280574
rect 178266 244658 178502 244894
rect 178586 244658 178822 244894
rect 178266 244338 178502 244574
rect 178586 244338 178822 244574
rect 178266 208658 178502 208894
rect 178586 208658 178822 208894
rect 178266 208338 178502 208574
rect 178586 208338 178822 208574
rect 178266 172658 178502 172894
rect 178586 172658 178822 172894
rect 178266 172338 178502 172574
rect 178586 172338 178822 172574
rect 178266 136658 178502 136894
rect 178586 136658 178822 136894
rect 178266 136338 178502 136574
rect 178586 136338 178822 136574
rect 178266 100658 178502 100894
rect 178586 100658 178822 100894
rect 178266 100338 178502 100574
rect 178586 100338 178822 100574
rect 178266 64658 178502 64894
rect 178586 64658 178822 64894
rect 178266 64338 178502 64574
rect 178586 64338 178822 64574
rect 178266 28658 178502 28894
rect 178586 28658 178822 28894
rect 178266 28338 178502 28574
rect 178586 28338 178822 28574
rect 180826 704602 181062 704838
rect 181146 704602 181382 704838
rect 180826 704282 181062 704518
rect 181146 704282 181382 704518
rect 180826 687218 181062 687454
rect 181146 687218 181382 687454
rect 180826 686898 181062 687134
rect 181146 686898 181382 687134
rect 180826 651218 181062 651454
rect 181146 651218 181382 651454
rect 180826 650898 181062 651134
rect 181146 650898 181382 651134
rect 180826 615218 181062 615454
rect 181146 615218 181382 615454
rect 180826 614898 181062 615134
rect 181146 614898 181382 615134
rect 180826 579218 181062 579454
rect 181146 579218 181382 579454
rect 180826 578898 181062 579134
rect 181146 578898 181382 579134
rect 180826 543218 181062 543454
rect 181146 543218 181382 543454
rect 180826 542898 181062 543134
rect 181146 542898 181382 543134
rect 180826 507218 181062 507454
rect 181146 507218 181382 507454
rect 180826 506898 181062 507134
rect 181146 506898 181382 507134
rect 180826 471218 181062 471454
rect 181146 471218 181382 471454
rect 180826 470898 181062 471134
rect 181146 470898 181382 471134
rect 180826 435218 181062 435454
rect 181146 435218 181382 435454
rect 180826 434898 181062 435134
rect 181146 434898 181382 435134
rect 180826 399218 181062 399454
rect 181146 399218 181382 399454
rect 180826 398898 181062 399134
rect 181146 398898 181382 399134
rect 180826 363218 181062 363454
rect 181146 363218 181382 363454
rect 180826 362898 181062 363134
rect 181146 362898 181382 363134
rect 180826 327218 181062 327454
rect 181146 327218 181382 327454
rect 180826 326898 181062 327134
rect 181146 326898 181382 327134
rect 180826 291218 181062 291454
rect 181146 291218 181382 291454
rect 180826 290898 181062 291134
rect 181146 290898 181382 291134
rect 180826 255218 181062 255454
rect 181146 255218 181382 255454
rect 180826 254898 181062 255134
rect 181146 254898 181382 255134
rect 180826 219218 181062 219454
rect 181146 219218 181382 219454
rect 180826 218898 181062 219134
rect 181146 218898 181382 219134
rect 180826 183218 181062 183454
rect 181146 183218 181382 183454
rect 180826 182898 181062 183134
rect 181146 182898 181382 183134
rect 180826 147218 181062 147454
rect 181146 147218 181382 147454
rect 180826 146898 181062 147134
rect 181146 146898 181382 147134
rect 180826 111218 181062 111454
rect 181146 111218 181382 111454
rect 180826 110898 181062 111134
rect 181146 110898 181382 111134
rect 180826 75218 181062 75454
rect 181146 75218 181382 75454
rect 180826 74898 181062 75134
rect 181146 74898 181382 75134
rect 180826 39218 181062 39454
rect 181146 39218 181382 39454
rect 180826 38898 181062 39134
rect 181146 38898 181382 39134
rect 180826 3218 181062 3454
rect 181146 3218 181382 3454
rect 180826 2898 181062 3134
rect 181146 2898 181382 3134
rect 180826 -582 181062 -346
rect 181146 -582 181382 -346
rect 180826 -902 181062 -666
rect 181146 -902 181382 -666
rect 191986 710362 192222 710598
rect 192306 710362 192542 710598
rect 191986 710042 192222 710278
rect 192306 710042 192542 710278
rect 188266 708442 188502 708678
rect 188586 708442 188822 708678
rect 188266 708122 188502 708358
rect 188586 708122 188822 708358
rect 181986 680378 182222 680614
rect 182306 680378 182542 680614
rect 181986 680058 182222 680294
rect 182306 680058 182542 680294
rect 181986 644378 182222 644614
rect 182306 644378 182542 644614
rect 181986 644058 182222 644294
rect 182306 644058 182542 644294
rect 181986 608378 182222 608614
rect 182306 608378 182542 608614
rect 181986 608058 182222 608294
rect 182306 608058 182542 608294
rect 181986 572378 182222 572614
rect 182306 572378 182542 572614
rect 181986 572058 182222 572294
rect 182306 572058 182542 572294
rect 181986 536378 182222 536614
rect 182306 536378 182542 536614
rect 181986 536058 182222 536294
rect 182306 536058 182542 536294
rect 181986 500378 182222 500614
rect 182306 500378 182542 500614
rect 181986 500058 182222 500294
rect 182306 500058 182542 500294
rect 181986 464378 182222 464614
rect 182306 464378 182542 464614
rect 181986 464058 182222 464294
rect 182306 464058 182542 464294
rect 181986 428378 182222 428614
rect 182306 428378 182542 428614
rect 181986 428058 182222 428294
rect 182306 428058 182542 428294
rect 181986 392378 182222 392614
rect 182306 392378 182542 392614
rect 181986 392058 182222 392294
rect 182306 392058 182542 392294
rect 181986 356378 182222 356614
rect 182306 356378 182542 356614
rect 181986 356058 182222 356294
rect 182306 356058 182542 356294
rect 181986 320378 182222 320614
rect 182306 320378 182542 320614
rect 181986 320058 182222 320294
rect 182306 320058 182542 320294
rect 181986 284378 182222 284614
rect 182306 284378 182542 284614
rect 181986 284058 182222 284294
rect 182306 284058 182542 284294
rect 181986 248378 182222 248614
rect 182306 248378 182542 248614
rect 181986 248058 182222 248294
rect 182306 248058 182542 248294
rect 181986 212378 182222 212614
rect 182306 212378 182542 212614
rect 181986 212058 182222 212294
rect 182306 212058 182542 212294
rect 181986 176378 182222 176614
rect 182306 176378 182542 176614
rect 181986 176058 182222 176294
rect 182306 176058 182542 176294
rect 181986 140378 182222 140614
rect 182306 140378 182542 140614
rect 181986 140058 182222 140294
rect 182306 140058 182542 140294
rect 181986 104378 182222 104614
rect 182306 104378 182542 104614
rect 181986 104058 182222 104294
rect 182306 104058 182542 104294
rect 181986 68378 182222 68614
rect 182306 68378 182542 68614
rect 181986 68058 182222 68294
rect 182306 68058 182542 68294
rect 181986 32378 182222 32614
rect 182306 32378 182542 32614
rect 181986 32058 182222 32294
rect 182306 32058 182542 32294
rect 178266 -5382 178502 -5146
rect 178586 -5382 178822 -5146
rect 178266 -5702 178502 -5466
rect 178586 -5702 178822 -5466
rect 171986 -6342 172222 -6106
rect 172306 -6342 172542 -6106
rect 171986 -6662 172222 -6426
rect 172306 -6662 172542 -6426
rect 184546 706522 184782 706758
rect 184866 706522 185102 706758
rect 184546 706202 184782 706438
rect 184866 706202 185102 706438
rect 184546 690938 184782 691174
rect 184866 690938 185102 691174
rect 184546 690618 184782 690854
rect 184866 690618 185102 690854
rect 184546 654938 184782 655174
rect 184866 654938 185102 655174
rect 184546 654618 184782 654854
rect 184866 654618 185102 654854
rect 184546 618938 184782 619174
rect 184866 618938 185102 619174
rect 184546 618618 184782 618854
rect 184866 618618 185102 618854
rect 184546 582938 184782 583174
rect 184866 582938 185102 583174
rect 184546 582618 184782 582854
rect 184866 582618 185102 582854
rect 184546 546938 184782 547174
rect 184866 546938 185102 547174
rect 184546 546618 184782 546854
rect 184866 546618 185102 546854
rect 184546 510938 184782 511174
rect 184866 510938 185102 511174
rect 184546 510618 184782 510854
rect 184866 510618 185102 510854
rect 184546 474938 184782 475174
rect 184866 474938 185102 475174
rect 184546 474618 184782 474854
rect 184866 474618 185102 474854
rect 184546 438938 184782 439174
rect 184866 438938 185102 439174
rect 184546 438618 184782 438854
rect 184866 438618 185102 438854
rect 184546 402938 184782 403174
rect 184866 402938 185102 403174
rect 184546 402618 184782 402854
rect 184866 402618 185102 402854
rect 184546 366938 184782 367174
rect 184866 366938 185102 367174
rect 184546 366618 184782 366854
rect 184866 366618 185102 366854
rect 184546 330938 184782 331174
rect 184866 330938 185102 331174
rect 184546 330618 184782 330854
rect 184866 330618 185102 330854
rect 184546 294938 184782 295174
rect 184866 294938 185102 295174
rect 184546 294618 184782 294854
rect 184866 294618 185102 294854
rect 184546 258938 184782 259174
rect 184866 258938 185102 259174
rect 184546 258618 184782 258854
rect 184866 258618 185102 258854
rect 184546 222938 184782 223174
rect 184866 222938 185102 223174
rect 184546 222618 184782 222854
rect 184866 222618 185102 222854
rect 184546 186938 184782 187174
rect 184866 186938 185102 187174
rect 184546 186618 184782 186854
rect 184866 186618 185102 186854
rect 184546 150938 184782 151174
rect 184866 150938 185102 151174
rect 184546 150618 184782 150854
rect 184866 150618 185102 150854
rect 184546 114938 184782 115174
rect 184866 114938 185102 115174
rect 184546 114618 184782 114854
rect 184866 114618 185102 114854
rect 184546 78938 184782 79174
rect 184866 78938 185102 79174
rect 184546 78618 184782 78854
rect 184866 78618 185102 78854
rect 184546 42938 184782 43174
rect 184866 42938 185102 43174
rect 184546 42618 184782 42854
rect 184866 42618 185102 42854
rect 184546 6938 184782 7174
rect 184866 6938 185102 7174
rect 184546 6618 184782 6854
rect 184866 6618 185102 6854
rect 184546 -2502 184782 -2266
rect 184866 -2502 185102 -2266
rect 184546 -2822 184782 -2586
rect 184866 -2822 185102 -2586
rect 188266 694658 188502 694894
rect 188586 694658 188822 694894
rect 188266 694338 188502 694574
rect 188586 694338 188822 694574
rect 188266 658658 188502 658894
rect 188586 658658 188822 658894
rect 188266 658338 188502 658574
rect 188586 658338 188822 658574
rect 188266 622658 188502 622894
rect 188586 622658 188822 622894
rect 188266 622338 188502 622574
rect 188586 622338 188822 622574
rect 188266 586658 188502 586894
rect 188586 586658 188822 586894
rect 188266 586338 188502 586574
rect 188586 586338 188822 586574
rect 188266 550658 188502 550894
rect 188586 550658 188822 550894
rect 188266 550338 188502 550574
rect 188586 550338 188822 550574
rect 188266 514658 188502 514894
rect 188586 514658 188822 514894
rect 188266 514338 188502 514574
rect 188586 514338 188822 514574
rect 188266 478658 188502 478894
rect 188586 478658 188822 478894
rect 188266 478338 188502 478574
rect 188586 478338 188822 478574
rect 188266 442658 188502 442894
rect 188586 442658 188822 442894
rect 188266 442338 188502 442574
rect 188586 442338 188822 442574
rect 188266 406658 188502 406894
rect 188586 406658 188822 406894
rect 188266 406338 188502 406574
rect 188586 406338 188822 406574
rect 188266 370658 188502 370894
rect 188586 370658 188822 370894
rect 188266 370338 188502 370574
rect 188586 370338 188822 370574
rect 188266 334658 188502 334894
rect 188586 334658 188822 334894
rect 188266 334338 188502 334574
rect 188586 334338 188822 334574
rect 188266 298658 188502 298894
rect 188586 298658 188822 298894
rect 188266 298338 188502 298574
rect 188586 298338 188822 298574
rect 188266 262658 188502 262894
rect 188586 262658 188822 262894
rect 188266 262338 188502 262574
rect 188586 262338 188822 262574
rect 188266 226658 188502 226894
rect 188586 226658 188822 226894
rect 188266 226338 188502 226574
rect 188586 226338 188822 226574
rect 188266 190658 188502 190894
rect 188586 190658 188822 190894
rect 188266 190338 188502 190574
rect 188586 190338 188822 190574
rect 188266 154658 188502 154894
rect 188586 154658 188822 154894
rect 188266 154338 188502 154574
rect 188586 154338 188822 154574
rect 188266 118658 188502 118894
rect 188586 118658 188822 118894
rect 188266 118338 188502 118574
rect 188586 118338 188822 118574
rect 188266 82658 188502 82894
rect 188586 82658 188822 82894
rect 188266 82338 188502 82574
rect 188586 82338 188822 82574
rect 188266 46658 188502 46894
rect 188586 46658 188822 46894
rect 188266 46338 188502 46574
rect 188586 46338 188822 46574
rect 188266 10658 188502 10894
rect 188586 10658 188822 10894
rect 188266 10338 188502 10574
rect 188586 10338 188822 10574
rect 190826 705562 191062 705798
rect 191146 705562 191382 705798
rect 190826 705242 191062 705478
rect 191146 705242 191382 705478
rect 190826 669218 191062 669454
rect 191146 669218 191382 669454
rect 190826 668898 191062 669134
rect 191146 668898 191382 669134
rect 190826 633218 191062 633454
rect 191146 633218 191382 633454
rect 190826 632898 191062 633134
rect 191146 632898 191382 633134
rect 190826 597218 191062 597454
rect 191146 597218 191382 597454
rect 190826 596898 191062 597134
rect 191146 596898 191382 597134
rect 190826 561218 191062 561454
rect 191146 561218 191382 561454
rect 190826 560898 191062 561134
rect 191146 560898 191382 561134
rect 190826 525218 191062 525454
rect 191146 525218 191382 525454
rect 190826 524898 191062 525134
rect 191146 524898 191382 525134
rect 190826 489218 191062 489454
rect 191146 489218 191382 489454
rect 190826 488898 191062 489134
rect 191146 488898 191382 489134
rect 190826 453218 191062 453454
rect 191146 453218 191382 453454
rect 190826 452898 191062 453134
rect 191146 452898 191382 453134
rect 190826 417218 191062 417454
rect 191146 417218 191382 417454
rect 190826 416898 191062 417134
rect 191146 416898 191382 417134
rect 190826 381218 191062 381454
rect 191146 381218 191382 381454
rect 190826 380898 191062 381134
rect 191146 380898 191382 381134
rect 190826 345218 191062 345454
rect 191146 345218 191382 345454
rect 190826 344898 191062 345134
rect 191146 344898 191382 345134
rect 190826 309218 191062 309454
rect 191146 309218 191382 309454
rect 190826 308898 191062 309134
rect 191146 308898 191382 309134
rect 190826 273218 191062 273454
rect 191146 273218 191382 273454
rect 190826 272898 191062 273134
rect 191146 272898 191382 273134
rect 190826 237218 191062 237454
rect 191146 237218 191382 237454
rect 190826 236898 191062 237134
rect 191146 236898 191382 237134
rect 190826 201218 191062 201454
rect 191146 201218 191382 201454
rect 190826 200898 191062 201134
rect 191146 200898 191382 201134
rect 190826 165218 191062 165454
rect 191146 165218 191382 165454
rect 190826 164898 191062 165134
rect 191146 164898 191382 165134
rect 190826 129218 191062 129454
rect 191146 129218 191382 129454
rect 190826 128898 191062 129134
rect 191146 128898 191382 129134
rect 190826 93218 191062 93454
rect 191146 93218 191382 93454
rect 190826 92898 191062 93134
rect 191146 92898 191382 93134
rect 190826 57218 191062 57454
rect 191146 57218 191382 57454
rect 190826 56898 191062 57134
rect 191146 56898 191382 57134
rect 190826 21218 191062 21454
rect 191146 21218 191382 21454
rect 190826 20898 191062 21134
rect 191146 20898 191382 21134
rect 190826 -1542 191062 -1306
rect 191146 -1542 191382 -1306
rect 190826 -1862 191062 -1626
rect 191146 -1862 191382 -1626
rect 201986 711322 202222 711558
rect 202306 711322 202542 711558
rect 201986 711002 202222 711238
rect 202306 711002 202542 711238
rect 198266 709402 198502 709638
rect 198586 709402 198822 709638
rect 198266 709082 198502 709318
rect 198586 709082 198822 709318
rect 191986 698378 192222 698614
rect 192306 698378 192542 698614
rect 191986 698058 192222 698294
rect 192306 698058 192542 698294
rect 191986 662378 192222 662614
rect 192306 662378 192542 662614
rect 191986 662058 192222 662294
rect 192306 662058 192542 662294
rect 191986 626378 192222 626614
rect 192306 626378 192542 626614
rect 191986 626058 192222 626294
rect 192306 626058 192542 626294
rect 191986 590378 192222 590614
rect 192306 590378 192542 590614
rect 191986 590058 192222 590294
rect 192306 590058 192542 590294
rect 191986 554378 192222 554614
rect 192306 554378 192542 554614
rect 191986 554058 192222 554294
rect 192306 554058 192542 554294
rect 191986 518378 192222 518614
rect 192306 518378 192542 518614
rect 191986 518058 192222 518294
rect 192306 518058 192542 518294
rect 191986 482378 192222 482614
rect 192306 482378 192542 482614
rect 191986 482058 192222 482294
rect 192306 482058 192542 482294
rect 191986 446378 192222 446614
rect 192306 446378 192542 446614
rect 191986 446058 192222 446294
rect 192306 446058 192542 446294
rect 191986 410378 192222 410614
rect 192306 410378 192542 410614
rect 191986 410058 192222 410294
rect 192306 410058 192542 410294
rect 191986 374378 192222 374614
rect 192306 374378 192542 374614
rect 191986 374058 192222 374294
rect 192306 374058 192542 374294
rect 191986 338378 192222 338614
rect 192306 338378 192542 338614
rect 191986 338058 192222 338294
rect 192306 338058 192542 338294
rect 191986 302378 192222 302614
rect 192306 302378 192542 302614
rect 191986 302058 192222 302294
rect 192306 302058 192542 302294
rect 191986 266378 192222 266614
rect 192306 266378 192542 266614
rect 191986 266058 192222 266294
rect 192306 266058 192542 266294
rect 191986 230378 192222 230614
rect 192306 230378 192542 230614
rect 191986 230058 192222 230294
rect 192306 230058 192542 230294
rect 191986 194378 192222 194614
rect 192306 194378 192542 194614
rect 191986 194058 192222 194294
rect 192306 194058 192542 194294
rect 191986 158378 192222 158614
rect 192306 158378 192542 158614
rect 191986 158058 192222 158294
rect 192306 158058 192542 158294
rect 191986 122378 192222 122614
rect 192306 122378 192542 122614
rect 191986 122058 192222 122294
rect 192306 122058 192542 122294
rect 191986 86378 192222 86614
rect 192306 86378 192542 86614
rect 191986 86058 192222 86294
rect 192306 86058 192542 86294
rect 191986 50378 192222 50614
rect 192306 50378 192542 50614
rect 191986 50058 192222 50294
rect 192306 50058 192542 50294
rect 191986 14378 192222 14614
rect 192306 14378 192542 14614
rect 191986 14058 192222 14294
rect 192306 14058 192542 14294
rect 188266 -4422 188502 -4186
rect 188586 -4422 188822 -4186
rect 188266 -4742 188502 -4506
rect 188586 -4742 188822 -4506
rect 181986 -7302 182222 -7066
rect 182306 -7302 182542 -7066
rect 181986 -7622 182222 -7386
rect 182306 -7622 182542 -7386
rect 194546 707482 194782 707718
rect 194866 707482 195102 707718
rect 194546 707162 194782 707398
rect 194866 707162 195102 707398
rect 194546 672938 194782 673174
rect 194866 672938 195102 673174
rect 194546 672618 194782 672854
rect 194866 672618 195102 672854
rect 194546 636938 194782 637174
rect 194866 636938 195102 637174
rect 194546 636618 194782 636854
rect 194866 636618 195102 636854
rect 194546 600938 194782 601174
rect 194866 600938 195102 601174
rect 194546 600618 194782 600854
rect 194866 600618 195102 600854
rect 194546 564938 194782 565174
rect 194866 564938 195102 565174
rect 194546 564618 194782 564854
rect 194866 564618 195102 564854
rect 194546 528938 194782 529174
rect 194866 528938 195102 529174
rect 194546 528618 194782 528854
rect 194866 528618 195102 528854
rect 194546 492938 194782 493174
rect 194866 492938 195102 493174
rect 194546 492618 194782 492854
rect 194866 492618 195102 492854
rect 194546 456938 194782 457174
rect 194866 456938 195102 457174
rect 194546 456618 194782 456854
rect 194866 456618 195102 456854
rect 194546 420938 194782 421174
rect 194866 420938 195102 421174
rect 194546 420618 194782 420854
rect 194866 420618 195102 420854
rect 194546 384938 194782 385174
rect 194866 384938 195102 385174
rect 194546 384618 194782 384854
rect 194866 384618 195102 384854
rect 194546 348938 194782 349174
rect 194866 348938 195102 349174
rect 194546 348618 194782 348854
rect 194866 348618 195102 348854
rect 194546 312938 194782 313174
rect 194866 312938 195102 313174
rect 194546 312618 194782 312854
rect 194866 312618 195102 312854
rect 194546 276938 194782 277174
rect 194866 276938 195102 277174
rect 194546 276618 194782 276854
rect 194866 276618 195102 276854
rect 194546 240938 194782 241174
rect 194866 240938 195102 241174
rect 194546 240618 194782 240854
rect 194866 240618 195102 240854
rect 194546 204938 194782 205174
rect 194866 204938 195102 205174
rect 194546 204618 194782 204854
rect 194866 204618 195102 204854
rect 194546 168938 194782 169174
rect 194866 168938 195102 169174
rect 194546 168618 194782 168854
rect 194866 168618 195102 168854
rect 194546 132938 194782 133174
rect 194866 132938 195102 133174
rect 194546 132618 194782 132854
rect 194866 132618 195102 132854
rect 194546 96938 194782 97174
rect 194866 96938 195102 97174
rect 194546 96618 194782 96854
rect 194866 96618 195102 96854
rect 194546 60938 194782 61174
rect 194866 60938 195102 61174
rect 194546 60618 194782 60854
rect 194866 60618 195102 60854
rect 194546 24938 194782 25174
rect 194866 24938 195102 25174
rect 194546 24618 194782 24854
rect 194866 24618 195102 24854
rect 194546 -3462 194782 -3226
rect 194866 -3462 195102 -3226
rect 194546 -3782 194782 -3546
rect 194866 -3782 195102 -3546
rect 198266 676658 198502 676894
rect 198586 676658 198822 676894
rect 198266 676338 198502 676574
rect 198586 676338 198822 676574
rect 198266 640658 198502 640894
rect 198586 640658 198822 640894
rect 198266 640338 198502 640574
rect 198586 640338 198822 640574
rect 198266 604658 198502 604894
rect 198586 604658 198822 604894
rect 198266 604338 198502 604574
rect 198586 604338 198822 604574
rect 198266 568658 198502 568894
rect 198586 568658 198822 568894
rect 198266 568338 198502 568574
rect 198586 568338 198822 568574
rect 198266 532658 198502 532894
rect 198586 532658 198822 532894
rect 198266 532338 198502 532574
rect 198586 532338 198822 532574
rect 198266 496658 198502 496894
rect 198586 496658 198822 496894
rect 198266 496338 198502 496574
rect 198586 496338 198822 496574
rect 198266 460658 198502 460894
rect 198586 460658 198822 460894
rect 198266 460338 198502 460574
rect 198586 460338 198822 460574
rect 198266 424658 198502 424894
rect 198586 424658 198822 424894
rect 198266 424338 198502 424574
rect 198586 424338 198822 424574
rect 198266 388658 198502 388894
rect 198586 388658 198822 388894
rect 198266 388338 198502 388574
rect 198586 388338 198822 388574
rect 198266 352658 198502 352894
rect 198586 352658 198822 352894
rect 198266 352338 198502 352574
rect 198586 352338 198822 352574
rect 198266 316658 198502 316894
rect 198586 316658 198822 316894
rect 198266 316338 198502 316574
rect 198586 316338 198822 316574
rect 198266 280658 198502 280894
rect 198586 280658 198822 280894
rect 198266 280338 198502 280574
rect 198586 280338 198822 280574
rect 198266 244658 198502 244894
rect 198586 244658 198822 244894
rect 198266 244338 198502 244574
rect 198586 244338 198822 244574
rect 198266 208658 198502 208894
rect 198586 208658 198822 208894
rect 198266 208338 198502 208574
rect 198586 208338 198822 208574
rect 198266 172658 198502 172894
rect 198586 172658 198822 172894
rect 198266 172338 198502 172574
rect 198586 172338 198822 172574
rect 198266 136658 198502 136894
rect 198586 136658 198822 136894
rect 198266 136338 198502 136574
rect 198586 136338 198822 136574
rect 198266 100658 198502 100894
rect 198586 100658 198822 100894
rect 198266 100338 198502 100574
rect 198586 100338 198822 100574
rect 198266 64658 198502 64894
rect 198586 64658 198822 64894
rect 198266 64338 198502 64574
rect 198586 64338 198822 64574
rect 198266 28658 198502 28894
rect 198586 28658 198822 28894
rect 198266 28338 198502 28574
rect 198586 28338 198822 28574
rect 200826 704602 201062 704838
rect 201146 704602 201382 704838
rect 200826 704282 201062 704518
rect 201146 704282 201382 704518
rect 200826 687218 201062 687454
rect 201146 687218 201382 687454
rect 200826 686898 201062 687134
rect 201146 686898 201382 687134
rect 200826 651218 201062 651454
rect 201146 651218 201382 651454
rect 200826 650898 201062 651134
rect 201146 650898 201382 651134
rect 200826 615218 201062 615454
rect 201146 615218 201382 615454
rect 200826 614898 201062 615134
rect 201146 614898 201382 615134
rect 200826 579218 201062 579454
rect 201146 579218 201382 579454
rect 200826 578898 201062 579134
rect 201146 578898 201382 579134
rect 200826 543218 201062 543454
rect 201146 543218 201382 543454
rect 200826 542898 201062 543134
rect 201146 542898 201382 543134
rect 200826 507218 201062 507454
rect 201146 507218 201382 507454
rect 200826 506898 201062 507134
rect 201146 506898 201382 507134
rect 200826 471218 201062 471454
rect 201146 471218 201382 471454
rect 200826 470898 201062 471134
rect 201146 470898 201382 471134
rect 200826 435218 201062 435454
rect 201146 435218 201382 435454
rect 200826 434898 201062 435134
rect 201146 434898 201382 435134
rect 200826 399218 201062 399454
rect 201146 399218 201382 399454
rect 200826 398898 201062 399134
rect 201146 398898 201382 399134
rect 200826 363218 201062 363454
rect 201146 363218 201382 363454
rect 200826 362898 201062 363134
rect 201146 362898 201382 363134
rect 200826 327218 201062 327454
rect 201146 327218 201382 327454
rect 200826 326898 201062 327134
rect 201146 326898 201382 327134
rect 200826 291218 201062 291454
rect 201146 291218 201382 291454
rect 200826 290898 201062 291134
rect 201146 290898 201382 291134
rect 200826 255218 201062 255454
rect 201146 255218 201382 255454
rect 200826 254898 201062 255134
rect 201146 254898 201382 255134
rect 200826 219218 201062 219454
rect 201146 219218 201382 219454
rect 200826 218898 201062 219134
rect 201146 218898 201382 219134
rect 200826 183218 201062 183454
rect 201146 183218 201382 183454
rect 200826 182898 201062 183134
rect 201146 182898 201382 183134
rect 200826 147218 201062 147454
rect 201146 147218 201382 147454
rect 200826 146898 201062 147134
rect 201146 146898 201382 147134
rect 200826 111218 201062 111454
rect 201146 111218 201382 111454
rect 200826 110898 201062 111134
rect 201146 110898 201382 111134
rect 200826 75218 201062 75454
rect 201146 75218 201382 75454
rect 200826 74898 201062 75134
rect 201146 74898 201382 75134
rect 200826 39218 201062 39454
rect 201146 39218 201382 39454
rect 200826 38898 201062 39134
rect 201146 38898 201382 39134
rect 200826 3218 201062 3454
rect 201146 3218 201382 3454
rect 200826 2898 201062 3134
rect 201146 2898 201382 3134
rect 200826 -582 201062 -346
rect 201146 -582 201382 -346
rect 200826 -902 201062 -666
rect 201146 -902 201382 -666
rect 211986 710362 212222 710598
rect 212306 710362 212542 710598
rect 211986 710042 212222 710278
rect 212306 710042 212542 710278
rect 208266 708442 208502 708678
rect 208586 708442 208822 708678
rect 208266 708122 208502 708358
rect 208586 708122 208822 708358
rect 201986 680378 202222 680614
rect 202306 680378 202542 680614
rect 201986 680058 202222 680294
rect 202306 680058 202542 680294
rect 201986 644378 202222 644614
rect 202306 644378 202542 644614
rect 201986 644058 202222 644294
rect 202306 644058 202542 644294
rect 201986 608378 202222 608614
rect 202306 608378 202542 608614
rect 201986 608058 202222 608294
rect 202306 608058 202542 608294
rect 201986 572378 202222 572614
rect 202306 572378 202542 572614
rect 201986 572058 202222 572294
rect 202306 572058 202542 572294
rect 201986 536378 202222 536614
rect 202306 536378 202542 536614
rect 201986 536058 202222 536294
rect 202306 536058 202542 536294
rect 201986 500378 202222 500614
rect 202306 500378 202542 500614
rect 201986 500058 202222 500294
rect 202306 500058 202542 500294
rect 201986 464378 202222 464614
rect 202306 464378 202542 464614
rect 201986 464058 202222 464294
rect 202306 464058 202542 464294
rect 201986 428378 202222 428614
rect 202306 428378 202542 428614
rect 201986 428058 202222 428294
rect 202306 428058 202542 428294
rect 201986 392378 202222 392614
rect 202306 392378 202542 392614
rect 201986 392058 202222 392294
rect 202306 392058 202542 392294
rect 201986 356378 202222 356614
rect 202306 356378 202542 356614
rect 201986 356058 202222 356294
rect 202306 356058 202542 356294
rect 201986 320378 202222 320614
rect 202306 320378 202542 320614
rect 201986 320058 202222 320294
rect 202306 320058 202542 320294
rect 201986 284378 202222 284614
rect 202306 284378 202542 284614
rect 201986 284058 202222 284294
rect 202306 284058 202542 284294
rect 201986 248378 202222 248614
rect 202306 248378 202542 248614
rect 201986 248058 202222 248294
rect 202306 248058 202542 248294
rect 201986 212378 202222 212614
rect 202306 212378 202542 212614
rect 201986 212058 202222 212294
rect 202306 212058 202542 212294
rect 201986 176378 202222 176614
rect 202306 176378 202542 176614
rect 201986 176058 202222 176294
rect 202306 176058 202542 176294
rect 201986 140378 202222 140614
rect 202306 140378 202542 140614
rect 201986 140058 202222 140294
rect 202306 140058 202542 140294
rect 201986 104378 202222 104614
rect 202306 104378 202542 104614
rect 201986 104058 202222 104294
rect 202306 104058 202542 104294
rect 201986 68378 202222 68614
rect 202306 68378 202542 68614
rect 201986 68058 202222 68294
rect 202306 68058 202542 68294
rect 201986 32378 202222 32614
rect 202306 32378 202542 32614
rect 201986 32058 202222 32294
rect 202306 32058 202542 32294
rect 198266 -5382 198502 -5146
rect 198586 -5382 198822 -5146
rect 198266 -5702 198502 -5466
rect 198586 -5702 198822 -5466
rect 191986 -6342 192222 -6106
rect 192306 -6342 192542 -6106
rect 191986 -6662 192222 -6426
rect 192306 -6662 192542 -6426
rect 204546 706522 204782 706758
rect 204866 706522 205102 706758
rect 204546 706202 204782 706438
rect 204866 706202 205102 706438
rect 204546 690938 204782 691174
rect 204866 690938 205102 691174
rect 204546 690618 204782 690854
rect 204866 690618 205102 690854
rect 204546 654938 204782 655174
rect 204866 654938 205102 655174
rect 204546 654618 204782 654854
rect 204866 654618 205102 654854
rect 204546 618938 204782 619174
rect 204866 618938 205102 619174
rect 204546 618618 204782 618854
rect 204866 618618 205102 618854
rect 204546 582938 204782 583174
rect 204866 582938 205102 583174
rect 204546 582618 204782 582854
rect 204866 582618 205102 582854
rect 204546 546938 204782 547174
rect 204866 546938 205102 547174
rect 204546 546618 204782 546854
rect 204866 546618 205102 546854
rect 204546 510938 204782 511174
rect 204866 510938 205102 511174
rect 204546 510618 204782 510854
rect 204866 510618 205102 510854
rect 204546 474938 204782 475174
rect 204866 474938 205102 475174
rect 204546 474618 204782 474854
rect 204866 474618 205102 474854
rect 204546 438938 204782 439174
rect 204866 438938 205102 439174
rect 204546 438618 204782 438854
rect 204866 438618 205102 438854
rect 204546 402938 204782 403174
rect 204866 402938 205102 403174
rect 204546 402618 204782 402854
rect 204866 402618 205102 402854
rect 204546 366938 204782 367174
rect 204866 366938 205102 367174
rect 204546 366618 204782 366854
rect 204866 366618 205102 366854
rect 204546 330938 204782 331174
rect 204866 330938 205102 331174
rect 204546 330618 204782 330854
rect 204866 330618 205102 330854
rect 204546 294938 204782 295174
rect 204866 294938 205102 295174
rect 204546 294618 204782 294854
rect 204866 294618 205102 294854
rect 204546 258938 204782 259174
rect 204866 258938 205102 259174
rect 204546 258618 204782 258854
rect 204866 258618 205102 258854
rect 204546 222938 204782 223174
rect 204866 222938 205102 223174
rect 204546 222618 204782 222854
rect 204866 222618 205102 222854
rect 204546 186938 204782 187174
rect 204866 186938 205102 187174
rect 204546 186618 204782 186854
rect 204866 186618 205102 186854
rect 204546 150938 204782 151174
rect 204866 150938 205102 151174
rect 204546 150618 204782 150854
rect 204866 150618 205102 150854
rect 204546 114938 204782 115174
rect 204866 114938 205102 115174
rect 204546 114618 204782 114854
rect 204866 114618 205102 114854
rect 204546 78938 204782 79174
rect 204866 78938 205102 79174
rect 204546 78618 204782 78854
rect 204866 78618 205102 78854
rect 204546 42938 204782 43174
rect 204866 42938 205102 43174
rect 204546 42618 204782 42854
rect 204866 42618 205102 42854
rect 204546 6938 204782 7174
rect 204866 6938 205102 7174
rect 204546 6618 204782 6854
rect 204866 6618 205102 6854
rect 204546 -2502 204782 -2266
rect 204866 -2502 205102 -2266
rect 204546 -2822 204782 -2586
rect 204866 -2822 205102 -2586
rect 208266 694658 208502 694894
rect 208586 694658 208822 694894
rect 208266 694338 208502 694574
rect 208586 694338 208822 694574
rect 208266 658658 208502 658894
rect 208586 658658 208822 658894
rect 208266 658338 208502 658574
rect 208586 658338 208822 658574
rect 208266 622658 208502 622894
rect 208586 622658 208822 622894
rect 208266 622338 208502 622574
rect 208586 622338 208822 622574
rect 208266 586658 208502 586894
rect 208586 586658 208822 586894
rect 208266 586338 208502 586574
rect 208586 586338 208822 586574
rect 208266 550658 208502 550894
rect 208586 550658 208822 550894
rect 208266 550338 208502 550574
rect 208586 550338 208822 550574
rect 208266 514658 208502 514894
rect 208586 514658 208822 514894
rect 208266 514338 208502 514574
rect 208586 514338 208822 514574
rect 208266 478658 208502 478894
rect 208586 478658 208822 478894
rect 208266 478338 208502 478574
rect 208586 478338 208822 478574
rect 208266 442658 208502 442894
rect 208586 442658 208822 442894
rect 208266 442338 208502 442574
rect 208586 442338 208822 442574
rect 208266 406658 208502 406894
rect 208586 406658 208822 406894
rect 208266 406338 208502 406574
rect 208586 406338 208822 406574
rect 208266 370658 208502 370894
rect 208586 370658 208822 370894
rect 208266 370338 208502 370574
rect 208586 370338 208822 370574
rect 208266 334658 208502 334894
rect 208586 334658 208822 334894
rect 208266 334338 208502 334574
rect 208586 334338 208822 334574
rect 208266 298658 208502 298894
rect 208586 298658 208822 298894
rect 208266 298338 208502 298574
rect 208586 298338 208822 298574
rect 208266 262658 208502 262894
rect 208586 262658 208822 262894
rect 208266 262338 208502 262574
rect 208586 262338 208822 262574
rect 208266 226658 208502 226894
rect 208586 226658 208822 226894
rect 208266 226338 208502 226574
rect 208586 226338 208822 226574
rect 208266 190658 208502 190894
rect 208586 190658 208822 190894
rect 208266 190338 208502 190574
rect 208586 190338 208822 190574
rect 208266 154658 208502 154894
rect 208586 154658 208822 154894
rect 208266 154338 208502 154574
rect 208586 154338 208822 154574
rect 208266 118658 208502 118894
rect 208586 118658 208822 118894
rect 208266 118338 208502 118574
rect 208586 118338 208822 118574
rect 208266 82658 208502 82894
rect 208586 82658 208822 82894
rect 208266 82338 208502 82574
rect 208586 82338 208822 82574
rect 208266 46658 208502 46894
rect 208586 46658 208822 46894
rect 208266 46338 208502 46574
rect 208586 46338 208822 46574
rect 208266 10658 208502 10894
rect 208586 10658 208822 10894
rect 208266 10338 208502 10574
rect 208586 10338 208822 10574
rect 210826 705562 211062 705798
rect 211146 705562 211382 705798
rect 210826 705242 211062 705478
rect 211146 705242 211382 705478
rect 210826 669218 211062 669454
rect 211146 669218 211382 669454
rect 210826 668898 211062 669134
rect 211146 668898 211382 669134
rect 210826 633218 211062 633454
rect 211146 633218 211382 633454
rect 210826 632898 211062 633134
rect 211146 632898 211382 633134
rect 210826 597218 211062 597454
rect 211146 597218 211382 597454
rect 210826 596898 211062 597134
rect 211146 596898 211382 597134
rect 210826 561218 211062 561454
rect 211146 561218 211382 561454
rect 210826 560898 211062 561134
rect 211146 560898 211382 561134
rect 210826 525218 211062 525454
rect 211146 525218 211382 525454
rect 210826 524898 211062 525134
rect 211146 524898 211382 525134
rect 210826 489218 211062 489454
rect 211146 489218 211382 489454
rect 210826 488898 211062 489134
rect 211146 488898 211382 489134
rect 210826 453218 211062 453454
rect 211146 453218 211382 453454
rect 210826 452898 211062 453134
rect 211146 452898 211382 453134
rect 210826 417218 211062 417454
rect 211146 417218 211382 417454
rect 210826 416898 211062 417134
rect 211146 416898 211382 417134
rect 210826 381218 211062 381454
rect 211146 381218 211382 381454
rect 210826 380898 211062 381134
rect 211146 380898 211382 381134
rect 210826 345218 211062 345454
rect 211146 345218 211382 345454
rect 210826 344898 211062 345134
rect 211146 344898 211382 345134
rect 210826 309218 211062 309454
rect 211146 309218 211382 309454
rect 210826 308898 211062 309134
rect 211146 308898 211382 309134
rect 210826 273218 211062 273454
rect 211146 273218 211382 273454
rect 210826 272898 211062 273134
rect 211146 272898 211382 273134
rect 210826 237218 211062 237454
rect 211146 237218 211382 237454
rect 210826 236898 211062 237134
rect 211146 236898 211382 237134
rect 210826 201218 211062 201454
rect 211146 201218 211382 201454
rect 210826 200898 211062 201134
rect 211146 200898 211382 201134
rect 210826 165218 211062 165454
rect 211146 165218 211382 165454
rect 210826 164898 211062 165134
rect 211146 164898 211382 165134
rect 210826 129218 211062 129454
rect 211146 129218 211382 129454
rect 210826 128898 211062 129134
rect 211146 128898 211382 129134
rect 210826 93218 211062 93454
rect 211146 93218 211382 93454
rect 210826 92898 211062 93134
rect 211146 92898 211382 93134
rect 210826 57218 211062 57454
rect 211146 57218 211382 57454
rect 210826 56898 211062 57134
rect 211146 56898 211382 57134
rect 210826 21218 211062 21454
rect 211146 21218 211382 21454
rect 210826 20898 211062 21134
rect 211146 20898 211382 21134
rect 210826 -1542 211062 -1306
rect 211146 -1542 211382 -1306
rect 210826 -1862 211062 -1626
rect 211146 -1862 211382 -1626
rect 221986 711322 222222 711558
rect 222306 711322 222542 711558
rect 221986 711002 222222 711238
rect 222306 711002 222542 711238
rect 218266 709402 218502 709638
rect 218586 709402 218822 709638
rect 218266 709082 218502 709318
rect 218586 709082 218822 709318
rect 211986 698378 212222 698614
rect 212306 698378 212542 698614
rect 211986 698058 212222 698294
rect 212306 698058 212542 698294
rect 211986 662378 212222 662614
rect 212306 662378 212542 662614
rect 211986 662058 212222 662294
rect 212306 662058 212542 662294
rect 211986 626378 212222 626614
rect 212306 626378 212542 626614
rect 211986 626058 212222 626294
rect 212306 626058 212542 626294
rect 211986 590378 212222 590614
rect 212306 590378 212542 590614
rect 211986 590058 212222 590294
rect 212306 590058 212542 590294
rect 211986 554378 212222 554614
rect 212306 554378 212542 554614
rect 211986 554058 212222 554294
rect 212306 554058 212542 554294
rect 211986 518378 212222 518614
rect 212306 518378 212542 518614
rect 211986 518058 212222 518294
rect 212306 518058 212542 518294
rect 211986 482378 212222 482614
rect 212306 482378 212542 482614
rect 211986 482058 212222 482294
rect 212306 482058 212542 482294
rect 211986 446378 212222 446614
rect 212306 446378 212542 446614
rect 211986 446058 212222 446294
rect 212306 446058 212542 446294
rect 211986 410378 212222 410614
rect 212306 410378 212542 410614
rect 211986 410058 212222 410294
rect 212306 410058 212542 410294
rect 211986 374378 212222 374614
rect 212306 374378 212542 374614
rect 211986 374058 212222 374294
rect 212306 374058 212542 374294
rect 211986 338378 212222 338614
rect 212306 338378 212542 338614
rect 211986 338058 212222 338294
rect 212306 338058 212542 338294
rect 211986 302378 212222 302614
rect 212306 302378 212542 302614
rect 211986 302058 212222 302294
rect 212306 302058 212542 302294
rect 211986 266378 212222 266614
rect 212306 266378 212542 266614
rect 211986 266058 212222 266294
rect 212306 266058 212542 266294
rect 211986 230378 212222 230614
rect 212306 230378 212542 230614
rect 211986 230058 212222 230294
rect 212306 230058 212542 230294
rect 211986 194378 212222 194614
rect 212306 194378 212542 194614
rect 211986 194058 212222 194294
rect 212306 194058 212542 194294
rect 211986 158378 212222 158614
rect 212306 158378 212542 158614
rect 211986 158058 212222 158294
rect 212306 158058 212542 158294
rect 211986 122378 212222 122614
rect 212306 122378 212542 122614
rect 211986 122058 212222 122294
rect 212306 122058 212542 122294
rect 211986 86378 212222 86614
rect 212306 86378 212542 86614
rect 211986 86058 212222 86294
rect 212306 86058 212542 86294
rect 211986 50378 212222 50614
rect 212306 50378 212542 50614
rect 211986 50058 212222 50294
rect 212306 50058 212542 50294
rect 211986 14378 212222 14614
rect 212306 14378 212542 14614
rect 211986 14058 212222 14294
rect 212306 14058 212542 14294
rect 208266 -4422 208502 -4186
rect 208586 -4422 208822 -4186
rect 208266 -4742 208502 -4506
rect 208586 -4742 208822 -4506
rect 201986 -7302 202222 -7066
rect 202306 -7302 202542 -7066
rect 201986 -7622 202222 -7386
rect 202306 -7622 202542 -7386
rect 214546 707482 214782 707718
rect 214866 707482 215102 707718
rect 214546 707162 214782 707398
rect 214866 707162 215102 707398
rect 214546 672938 214782 673174
rect 214866 672938 215102 673174
rect 214546 672618 214782 672854
rect 214866 672618 215102 672854
rect 214546 636938 214782 637174
rect 214866 636938 215102 637174
rect 214546 636618 214782 636854
rect 214866 636618 215102 636854
rect 214546 600938 214782 601174
rect 214866 600938 215102 601174
rect 214546 600618 214782 600854
rect 214866 600618 215102 600854
rect 214546 564938 214782 565174
rect 214866 564938 215102 565174
rect 214546 564618 214782 564854
rect 214866 564618 215102 564854
rect 214546 528938 214782 529174
rect 214866 528938 215102 529174
rect 214546 528618 214782 528854
rect 214866 528618 215102 528854
rect 214546 492938 214782 493174
rect 214866 492938 215102 493174
rect 214546 492618 214782 492854
rect 214866 492618 215102 492854
rect 214546 456938 214782 457174
rect 214866 456938 215102 457174
rect 214546 456618 214782 456854
rect 214866 456618 215102 456854
rect 214546 420938 214782 421174
rect 214866 420938 215102 421174
rect 214546 420618 214782 420854
rect 214866 420618 215102 420854
rect 214546 384938 214782 385174
rect 214866 384938 215102 385174
rect 214546 384618 214782 384854
rect 214866 384618 215102 384854
rect 214546 348938 214782 349174
rect 214866 348938 215102 349174
rect 214546 348618 214782 348854
rect 214866 348618 215102 348854
rect 214546 312938 214782 313174
rect 214866 312938 215102 313174
rect 214546 312618 214782 312854
rect 214866 312618 215102 312854
rect 214546 276938 214782 277174
rect 214866 276938 215102 277174
rect 214546 276618 214782 276854
rect 214866 276618 215102 276854
rect 214546 240938 214782 241174
rect 214866 240938 215102 241174
rect 214546 240618 214782 240854
rect 214866 240618 215102 240854
rect 214546 204938 214782 205174
rect 214866 204938 215102 205174
rect 214546 204618 214782 204854
rect 214866 204618 215102 204854
rect 214546 168938 214782 169174
rect 214866 168938 215102 169174
rect 214546 168618 214782 168854
rect 214866 168618 215102 168854
rect 214546 132938 214782 133174
rect 214866 132938 215102 133174
rect 214546 132618 214782 132854
rect 214866 132618 215102 132854
rect 214546 96938 214782 97174
rect 214866 96938 215102 97174
rect 214546 96618 214782 96854
rect 214866 96618 215102 96854
rect 214546 60938 214782 61174
rect 214866 60938 215102 61174
rect 214546 60618 214782 60854
rect 214866 60618 215102 60854
rect 214546 24938 214782 25174
rect 214866 24938 215102 25174
rect 214546 24618 214782 24854
rect 214866 24618 215102 24854
rect 214546 -3462 214782 -3226
rect 214866 -3462 215102 -3226
rect 214546 -3782 214782 -3546
rect 214866 -3782 215102 -3546
rect 218266 676658 218502 676894
rect 218586 676658 218822 676894
rect 218266 676338 218502 676574
rect 218586 676338 218822 676574
rect 218266 640658 218502 640894
rect 218586 640658 218822 640894
rect 218266 640338 218502 640574
rect 218586 640338 218822 640574
rect 218266 604658 218502 604894
rect 218586 604658 218822 604894
rect 218266 604338 218502 604574
rect 218586 604338 218822 604574
rect 218266 568658 218502 568894
rect 218586 568658 218822 568894
rect 218266 568338 218502 568574
rect 218586 568338 218822 568574
rect 218266 532658 218502 532894
rect 218586 532658 218822 532894
rect 218266 532338 218502 532574
rect 218586 532338 218822 532574
rect 218266 496658 218502 496894
rect 218586 496658 218822 496894
rect 218266 496338 218502 496574
rect 218586 496338 218822 496574
rect 218266 460658 218502 460894
rect 218586 460658 218822 460894
rect 218266 460338 218502 460574
rect 218586 460338 218822 460574
rect 218266 424658 218502 424894
rect 218586 424658 218822 424894
rect 218266 424338 218502 424574
rect 218586 424338 218822 424574
rect 218266 388658 218502 388894
rect 218586 388658 218822 388894
rect 218266 388338 218502 388574
rect 218586 388338 218822 388574
rect 218266 352658 218502 352894
rect 218586 352658 218822 352894
rect 218266 352338 218502 352574
rect 218586 352338 218822 352574
rect 218266 316658 218502 316894
rect 218586 316658 218822 316894
rect 218266 316338 218502 316574
rect 218586 316338 218822 316574
rect 218266 280658 218502 280894
rect 218586 280658 218822 280894
rect 218266 280338 218502 280574
rect 218586 280338 218822 280574
rect 218266 244658 218502 244894
rect 218586 244658 218822 244894
rect 218266 244338 218502 244574
rect 218586 244338 218822 244574
rect 218266 208658 218502 208894
rect 218586 208658 218822 208894
rect 218266 208338 218502 208574
rect 218586 208338 218822 208574
rect 218266 172658 218502 172894
rect 218586 172658 218822 172894
rect 218266 172338 218502 172574
rect 218586 172338 218822 172574
rect 218266 136658 218502 136894
rect 218586 136658 218822 136894
rect 218266 136338 218502 136574
rect 218586 136338 218822 136574
rect 218266 100658 218502 100894
rect 218586 100658 218822 100894
rect 218266 100338 218502 100574
rect 218586 100338 218822 100574
rect 218266 64658 218502 64894
rect 218586 64658 218822 64894
rect 218266 64338 218502 64574
rect 218586 64338 218822 64574
rect 218266 28658 218502 28894
rect 218586 28658 218822 28894
rect 218266 28338 218502 28574
rect 218586 28338 218822 28574
rect 220826 704602 221062 704838
rect 221146 704602 221382 704838
rect 220826 704282 221062 704518
rect 221146 704282 221382 704518
rect 220826 687218 221062 687454
rect 221146 687218 221382 687454
rect 220826 686898 221062 687134
rect 221146 686898 221382 687134
rect 220826 651218 221062 651454
rect 221146 651218 221382 651454
rect 220826 650898 221062 651134
rect 221146 650898 221382 651134
rect 220826 615218 221062 615454
rect 221146 615218 221382 615454
rect 220826 614898 221062 615134
rect 221146 614898 221382 615134
rect 220826 579218 221062 579454
rect 221146 579218 221382 579454
rect 220826 578898 221062 579134
rect 221146 578898 221382 579134
rect 220826 543218 221062 543454
rect 221146 543218 221382 543454
rect 220826 542898 221062 543134
rect 221146 542898 221382 543134
rect 220826 507218 221062 507454
rect 221146 507218 221382 507454
rect 220826 506898 221062 507134
rect 221146 506898 221382 507134
rect 220826 471218 221062 471454
rect 221146 471218 221382 471454
rect 220826 470898 221062 471134
rect 221146 470898 221382 471134
rect 220826 435218 221062 435454
rect 221146 435218 221382 435454
rect 220826 434898 221062 435134
rect 221146 434898 221382 435134
rect 220826 399218 221062 399454
rect 221146 399218 221382 399454
rect 220826 398898 221062 399134
rect 221146 398898 221382 399134
rect 220826 363218 221062 363454
rect 221146 363218 221382 363454
rect 220826 362898 221062 363134
rect 221146 362898 221382 363134
rect 220826 327218 221062 327454
rect 221146 327218 221382 327454
rect 220826 326898 221062 327134
rect 221146 326898 221382 327134
rect 220826 291218 221062 291454
rect 221146 291218 221382 291454
rect 220826 290898 221062 291134
rect 221146 290898 221382 291134
rect 220826 255218 221062 255454
rect 221146 255218 221382 255454
rect 220826 254898 221062 255134
rect 221146 254898 221382 255134
rect 220826 219218 221062 219454
rect 221146 219218 221382 219454
rect 220826 218898 221062 219134
rect 221146 218898 221382 219134
rect 220826 183218 221062 183454
rect 221146 183218 221382 183454
rect 220826 182898 221062 183134
rect 221146 182898 221382 183134
rect 220826 147218 221062 147454
rect 221146 147218 221382 147454
rect 220826 146898 221062 147134
rect 221146 146898 221382 147134
rect 220826 111218 221062 111454
rect 221146 111218 221382 111454
rect 220826 110898 221062 111134
rect 221146 110898 221382 111134
rect 220826 75218 221062 75454
rect 221146 75218 221382 75454
rect 220826 74898 221062 75134
rect 221146 74898 221382 75134
rect 220826 39218 221062 39454
rect 221146 39218 221382 39454
rect 220826 38898 221062 39134
rect 221146 38898 221382 39134
rect 220826 3218 221062 3454
rect 221146 3218 221382 3454
rect 220826 2898 221062 3134
rect 221146 2898 221382 3134
rect 220826 -582 221062 -346
rect 221146 -582 221382 -346
rect 220826 -902 221062 -666
rect 221146 -902 221382 -666
rect 231986 710362 232222 710598
rect 232306 710362 232542 710598
rect 231986 710042 232222 710278
rect 232306 710042 232542 710278
rect 228266 708442 228502 708678
rect 228586 708442 228822 708678
rect 228266 708122 228502 708358
rect 228586 708122 228822 708358
rect 221986 680378 222222 680614
rect 222306 680378 222542 680614
rect 221986 680058 222222 680294
rect 222306 680058 222542 680294
rect 221986 644378 222222 644614
rect 222306 644378 222542 644614
rect 221986 644058 222222 644294
rect 222306 644058 222542 644294
rect 221986 608378 222222 608614
rect 222306 608378 222542 608614
rect 221986 608058 222222 608294
rect 222306 608058 222542 608294
rect 221986 572378 222222 572614
rect 222306 572378 222542 572614
rect 221986 572058 222222 572294
rect 222306 572058 222542 572294
rect 221986 536378 222222 536614
rect 222306 536378 222542 536614
rect 221986 536058 222222 536294
rect 222306 536058 222542 536294
rect 221986 500378 222222 500614
rect 222306 500378 222542 500614
rect 221986 500058 222222 500294
rect 222306 500058 222542 500294
rect 221986 464378 222222 464614
rect 222306 464378 222542 464614
rect 221986 464058 222222 464294
rect 222306 464058 222542 464294
rect 221986 428378 222222 428614
rect 222306 428378 222542 428614
rect 221986 428058 222222 428294
rect 222306 428058 222542 428294
rect 221986 392378 222222 392614
rect 222306 392378 222542 392614
rect 221986 392058 222222 392294
rect 222306 392058 222542 392294
rect 221986 356378 222222 356614
rect 222306 356378 222542 356614
rect 221986 356058 222222 356294
rect 222306 356058 222542 356294
rect 221986 320378 222222 320614
rect 222306 320378 222542 320614
rect 221986 320058 222222 320294
rect 222306 320058 222542 320294
rect 221986 284378 222222 284614
rect 222306 284378 222542 284614
rect 221986 284058 222222 284294
rect 222306 284058 222542 284294
rect 221986 248378 222222 248614
rect 222306 248378 222542 248614
rect 221986 248058 222222 248294
rect 222306 248058 222542 248294
rect 221986 212378 222222 212614
rect 222306 212378 222542 212614
rect 221986 212058 222222 212294
rect 222306 212058 222542 212294
rect 221986 176378 222222 176614
rect 222306 176378 222542 176614
rect 221986 176058 222222 176294
rect 222306 176058 222542 176294
rect 221986 140378 222222 140614
rect 222306 140378 222542 140614
rect 221986 140058 222222 140294
rect 222306 140058 222542 140294
rect 221986 104378 222222 104614
rect 222306 104378 222542 104614
rect 221986 104058 222222 104294
rect 222306 104058 222542 104294
rect 221986 68378 222222 68614
rect 222306 68378 222542 68614
rect 221986 68058 222222 68294
rect 222306 68058 222542 68294
rect 221986 32378 222222 32614
rect 222306 32378 222542 32614
rect 221986 32058 222222 32294
rect 222306 32058 222542 32294
rect 218266 -5382 218502 -5146
rect 218586 -5382 218822 -5146
rect 218266 -5702 218502 -5466
rect 218586 -5702 218822 -5466
rect 211986 -6342 212222 -6106
rect 212306 -6342 212542 -6106
rect 211986 -6662 212222 -6426
rect 212306 -6662 212542 -6426
rect 224546 706522 224782 706758
rect 224866 706522 225102 706758
rect 224546 706202 224782 706438
rect 224866 706202 225102 706438
rect 224546 690938 224782 691174
rect 224866 690938 225102 691174
rect 224546 690618 224782 690854
rect 224866 690618 225102 690854
rect 224546 654938 224782 655174
rect 224866 654938 225102 655174
rect 224546 654618 224782 654854
rect 224866 654618 225102 654854
rect 224546 618938 224782 619174
rect 224866 618938 225102 619174
rect 224546 618618 224782 618854
rect 224866 618618 225102 618854
rect 224546 582938 224782 583174
rect 224866 582938 225102 583174
rect 224546 582618 224782 582854
rect 224866 582618 225102 582854
rect 224546 546938 224782 547174
rect 224866 546938 225102 547174
rect 224546 546618 224782 546854
rect 224866 546618 225102 546854
rect 224546 510938 224782 511174
rect 224866 510938 225102 511174
rect 224546 510618 224782 510854
rect 224866 510618 225102 510854
rect 224546 474938 224782 475174
rect 224866 474938 225102 475174
rect 224546 474618 224782 474854
rect 224866 474618 225102 474854
rect 224546 438938 224782 439174
rect 224866 438938 225102 439174
rect 224546 438618 224782 438854
rect 224866 438618 225102 438854
rect 224546 402938 224782 403174
rect 224866 402938 225102 403174
rect 224546 402618 224782 402854
rect 224866 402618 225102 402854
rect 224546 366938 224782 367174
rect 224866 366938 225102 367174
rect 224546 366618 224782 366854
rect 224866 366618 225102 366854
rect 224546 330938 224782 331174
rect 224866 330938 225102 331174
rect 224546 330618 224782 330854
rect 224866 330618 225102 330854
rect 224546 294938 224782 295174
rect 224866 294938 225102 295174
rect 224546 294618 224782 294854
rect 224866 294618 225102 294854
rect 224546 258938 224782 259174
rect 224866 258938 225102 259174
rect 224546 258618 224782 258854
rect 224866 258618 225102 258854
rect 224546 222938 224782 223174
rect 224866 222938 225102 223174
rect 224546 222618 224782 222854
rect 224866 222618 225102 222854
rect 224546 186938 224782 187174
rect 224866 186938 225102 187174
rect 224546 186618 224782 186854
rect 224866 186618 225102 186854
rect 224546 150938 224782 151174
rect 224866 150938 225102 151174
rect 224546 150618 224782 150854
rect 224866 150618 225102 150854
rect 224546 114938 224782 115174
rect 224866 114938 225102 115174
rect 224546 114618 224782 114854
rect 224866 114618 225102 114854
rect 224546 78938 224782 79174
rect 224866 78938 225102 79174
rect 224546 78618 224782 78854
rect 224866 78618 225102 78854
rect 224546 42938 224782 43174
rect 224866 42938 225102 43174
rect 224546 42618 224782 42854
rect 224866 42618 225102 42854
rect 224546 6938 224782 7174
rect 224866 6938 225102 7174
rect 224546 6618 224782 6854
rect 224866 6618 225102 6854
rect 224546 -2502 224782 -2266
rect 224866 -2502 225102 -2266
rect 224546 -2822 224782 -2586
rect 224866 -2822 225102 -2586
rect 228266 694658 228502 694894
rect 228586 694658 228822 694894
rect 228266 694338 228502 694574
rect 228586 694338 228822 694574
rect 228266 658658 228502 658894
rect 228586 658658 228822 658894
rect 228266 658338 228502 658574
rect 228586 658338 228822 658574
rect 228266 622658 228502 622894
rect 228586 622658 228822 622894
rect 228266 622338 228502 622574
rect 228586 622338 228822 622574
rect 228266 586658 228502 586894
rect 228586 586658 228822 586894
rect 228266 586338 228502 586574
rect 228586 586338 228822 586574
rect 228266 550658 228502 550894
rect 228586 550658 228822 550894
rect 228266 550338 228502 550574
rect 228586 550338 228822 550574
rect 228266 514658 228502 514894
rect 228586 514658 228822 514894
rect 228266 514338 228502 514574
rect 228586 514338 228822 514574
rect 228266 478658 228502 478894
rect 228586 478658 228822 478894
rect 228266 478338 228502 478574
rect 228586 478338 228822 478574
rect 228266 442658 228502 442894
rect 228586 442658 228822 442894
rect 228266 442338 228502 442574
rect 228586 442338 228822 442574
rect 228266 406658 228502 406894
rect 228586 406658 228822 406894
rect 228266 406338 228502 406574
rect 228586 406338 228822 406574
rect 228266 370658 228502 370894
rect 228586 370658 228822 370894
rect 228266 370338 228502 370574
rect 228586 370338 228822 370574
rect 228266 334658 228502 334894
rect 228586 334658 228822 334894
rect 228266 334338 228502 334574
rect 228586 334338 228822 334574
rect 228266 298658 228502 298894
rect 228586 298658 228822 298894
rect 228266 298338 228502 298574
rect 228586 298338 228822 298574
rect 228266 262658 228502 262894
rect 228586 262658 228822 262894
rect 228266 262338 228502 262574
rect 228586 262338 228822 262574
rect 228266 226658 228502 226894
rect 228586 226658 228822 226894
rect 228266 226338 228502 226574
rect 228586 226338 228822 226574
rect 228266 190658 228502 190894
rect 228586 190658 228822 190894
rect 228266 190338 228502 190574
rect 228586 190338 228822 190574
rect 228266 154658 228502 154894
rect 228586 154658 228822 154894
rect 228266 154338 228502 154574
rect 228586 154338 228822 154574
rect 228266 118658 228502 118894
rect 228586 118658 228822 118894
rect 228266 118338 228502 118574
rect 228586 118338 228822 118574
rect 228266 82658 228502 82894
rect 228586 82658 228822 82894
rect 228266 82338 228502 82574
rect 228586 82338 228822 82574
rect 228266 46658 228502 46894
rect 228586 46658 228822 46894
rect 228266 46338 228502 46574
rect 228586 46338 228822 46574
rect 228266 10658 228502 10894
rect 228586 10658 228822 10894
rect 228266 10338 228502 10574
rect 228586 10338 228822 10574
rect 230826 705562 231062 705798
rect 231146 705562 231382 705798
rect 230826 705242 231062 705478
rect 231146 705242 231382 705478
rect 230826 669218 231062 669454
rect 231146 669218 231382 669454
rect 230826 668898 231062 669134
rect 231146 668898 231382 669134
rect 230826 633218 231062 633454
rect 231146 633218 231382 633454
rect 230826 632898 231062 633134
rect 231146 632898 231382 633134
rect 230826 597218 231062 597454
rect 231146 597218 231382 597454
rect 230826 596898 231062 597134
rect 231146 596898 231382 597134
rect 230826 561218 231062 561454
rect 231146 561218 231382 561454
rect 230826 560898 231062 561134
rect 231146 560898 231382 561134
rect 230826 525218 231062 525454
rect 231146 525218 231382 525454
rect 230826 524898 231062 525134
rect 231146 524898 231382 525134
rect 230826 489218 231062 489454
rect 231146 489218 231382 489454
rect 230826 488898 231062 489134
rect 231146 488898 231382 489134
rect 230826 453218 231062 453454
rect 231146 453218 231382 453454
rect 230826 452898 231062 453134
rect 231146 452898 231382 453134
rect 230826 417218 231062 417454
rect 231146 417218 231382 417454
rect 230826 416898 231062 417134
rect 231146 416898 231382 417134
rect 230826 381218 231062 381454
rect 231146 381218 231382 381454
rect 230826 380898 231062 381134
rect 231146 380898 231382 381134
rect 230826 345218 231062 345454
rect 231146 345218 231382 345454
rect 230826 344898 231062 345134
rect 231146 344898 231382 345134
rect 230826 309218 231062 309454
rect 231146 309218 231382 309454
rect 230826 308898 231062 309134
rect 231146 308898 231382 309134
rect 230826 273218 231062 273454
rect 231146 273218 231382 273454
rect 230826 272898 231062 273134
rect 231146 272898 231382 273134
rect 230826 237218 231062 237454
rect 231146 237218 231382 237454
rect 230826 236898 231062 237134
rect 231146 236898 231382 237134
rect 230826 201218 231062 201454
rect 231146 201218 231382 201454
rect 230826 200898 231062 201134
rect 231146 200898 231382 201134
rect 230826 165218 231062 165454
rect 231146 165218 231382 165454
rect 230826 164898 231062 165134
rect 231146 164898 231382 165134
rect 230826 129218 231062 129454
rect 231146 129218 231382 129454
rect 230826 128898 231062 129134
rect 231146 128898 231382 129134
rect 230826 93218 231062 93454
rect 231146 93218 231382 93454
rect 230826 92898 231062 93134
rect 231146 92898 231382 93134
rect 230826 57218 231062 57454
rect 231146 57218 231382 57454
rect 230826 56898 231062 57134
rect 231146 56898 231382 57134
rect 230826 21218 231062 21454
rect 231146 21218 231382 21454
rect 230826 20898 231062 21134
rect 231146 20898 231382 21134
rect 230826 -1542 231062 -1306
rect 231146 -1542 231382 -1306
rect 230826 -1862 231062 -1626
rect 231146 -1862 231382 -1626
rect 241986 711322 242222 711558
rect 242306 711322 242542 711558
rect 241986 711002 242222 711238
rect 242306 711002 242542 711238
rect 238266 709402 238502 709638
rect 238586 709402 238822 709638
rect 238266 709082 238502 709318
rect 238586 709082 238822 709318
rect 231986 698378 232222 698614
rect 232306 698378 232542 698614
rect 231986 698058 232222 698294
rect 232306 698058 232542 698294
rect 231986 662378 232222 662614
rect 232306 662378 232542 662614
rect 231986 662058 232222 662294
rect 232306 662058 232542 662294
rect 231986 626378 232222 626614
rect 232306 626378 232542 626614
rect 231986 626058 232222 626294
rect 232306 626058 232542 626294
rect 231986 590378 232222 590614
rect 232306 590378 232542 590614
rect 231986 590058 232222 590294
rect 232306 590058 232542 590294
rect 231986 554378 232222 554614
rect 232306 554378 232542 554614
rect 231986 554058 232222 554294
rect 232306 554058 232542 554294
rect 231986 518378 232222 518614
rect 232306 518378 232542 518614
rect 231986 518058 232222 518294
rect 232306 518058 232542 518294
rect 231986 482378 232222 482614
rect 232306 482378 232542 482614
rect 231986 482058 232222 482294
rect 232306 482058 232542 482294
rect 231986 446378 232222 446614
rect 232306 446378 232542 446614
rect 231986 446058 232222 446294
rect 232306 446058 232542 446294
rect 231986 410378 232222 410614
rect 232306 410378 232542 410614
rect 231986 410058 232222 410294
rect 232306 410058 232542 410294
rect 231986 374378 232222 374614
rect 232306 374378 232542 374614
rect 231986 374058 232222 374294
rect 232306 374058 232542 374294
rect 231986 338378 232222 338614
rect 232306 338378 232542 338614
rect 231986 338058 232222 338294
rect 232306 338058 232542 338294
rect 231986 302378 232222 302614
rect 232306 302378 232542 302614
rect 231986 302058 232222 302294
rect 232306 302058 232542 302294
rect 231986 266378 232222 266614
rect 232306 266378 232542 266614
rect 231986 266058 232222 266294
rect 232306 266058 232542 266294
rect 231986 230378 232222 230614
rect 232306 230378 232542 230614
rect 231986 230058 232222 230294
rect 232306 230058 232542 230294
rect 231986 194378 232222 194614
rect 232306 194378 232542 194614
rect 231986 194058 232222 194294
rect 232306 194058 232542 194294
rect 231986 158378 232222 158614
rect 232306 158378 232542 158614
rect 231986 158058 232222 158294
rect 232306 158058 232542 158294
rect 231986 122378 232222 122614
rect 232306 122378 232542 122614
rect 231986 122058 232222 122294
rect 232306 122058 232542 122294
rect 231986 86378 232222 86614
rect 232306 86378 232542 86614
rect 231986 86058 232222 86294
rect 232306 86058 232542 86294
rect 231986 50378 232222 50614
rect 232306 50378 232542 50614
rect 231986 50058 232222 50294
rect 232306 50058 232542 50294
rect 231986 14378 232222 14614
rect 232306 14378 232542 14614
rect 231986 14058 232222 14294
rect 232306 14058 232542 14294
rect 228266 -4422 228502 -4186
rect 228586 -4422 228822 -4186
rect 228266 -4742 228502 -4506
rect 228586 -4742 228822 -4506
rect 221986 -7302 222222 -7066
rect 222306 -7302 222542 -7066
rect 221986 -7622 222222 -7386
rect 222306 -7622 222542 -7386
rect 234546 707482 234782 707718
rect 234866 707482 235102 707718
rect 234546 707162 234782 707398
rect 234866 707162 235102 707398
rect 234546 672938 234782 673174
rect 234866 672938 235102 673174
rect 234546 672618 234782 672854
rect 234866 672618 235102 672854
rect 234546 636938 234782 637174
rect 234866 636938 235102 637174
rect 234546 636618 234782 636854
rect 234866 636618 235102 636854
rect 234546 600938 234782 601174
rect 234866 600938 235102 601174
rect 234546 600618 234782 600854
rect 234866 600618 235102 600854
rect 234546 564938 234782 565174
rect 234866 564938 235102 565174
rect 234546 564618 234782 564854
rect 234866 564618 235102 564854
rect 234546 528938 234782 529174
rect 234866 528938 235102 529174
rect 234546 528618 234782 528854
rect 234866 528618 235102 528854
rect 234546 492938 234782 493174
rect 234866 492938 235102 493174
rect 234546 492618 234782 492854
rect 234866 492618 235102 492854
rect 234546 456938 234782 457174
rect 234866 456938 235102 457174
rect 234546 456618 234782 456854
rect 234866 456618 235102 456854
rect 234546 420938 234782 421174
rect 234866 420938 235102 421174
rect 234546 420618 234782 420854
rect 234866 420618 235102 420854
rect 234546 384938 234782 385174
rect 234866 384938 235102 385174
rect 234546 384618 234782 384854
rect 234866 384618 235102 384854
rect 234546 348938 234782 349174
rect 234866 348938 235102 349174
rect 234546 348618 234782 348854
rect 234866 348618 235102 348854
rect 234546 312938 234782 313174
rect 234866 312938 235102 313174
rect 234546 312618 234782 312854
rect 234866 312618 235102 312854
rect 234546 276938 234782 277174
rect 234866 276938 235102 277174
rect 234546 276618 234782 276854
rect 234866 276618 235102 276854
rect 234546 240938 234782 241174
rect 234866 240938 235102 241174
rect 234546 240618 234782 240854
rect 234866 240618 235102 240854
rect 234546 204938 234782 205174
rect 234866 204938 235102 205174
rect 234546 204618 234782 204854
rect 234866 204618 235102 204854
rect 234546 168938 234782 169174
rect 234866 168938 235102 169174
rect 234546 168618 234782 168854
rect 234866 168618 235102 168854
rect 234546 132938 234782 133174
rect 234866 132938 235102 133174
rect 234546 132618 234782 132854
rect 234866 132618 235102 132854
rect 234546 96938 234782 97174
rect 234866 96938 235102 97174
rect 234546 96618 234782 96854
rect 234866 96618 235102 96854
rect 234546 60938 234782 61174
rect 234866 60938 235102 61174
rect 234546 60618 234782 60854
rect 234866 60618 235102 60854
rect 234546 24938 234782 25174
rect 234866 24938 235102 25174
rect 234546 24618 234782 24854
rect 234866 24618 235102 24854
rect 234546 -3462 234782 -3226
rect 234866 -3462 235102 -3226
rect 234546 -3782 234782 -3546
rect 234866 -3782 235102 -3546
rect 238266 676658 238502 676894
rect 238586 676658 238822 676894
rect 238266 676338 238502 676574
rect 238586 676338 238822 676574
rect 238266 640658 238502 640894
rect 238586 640658 238822 640894
rect 238266 640338 238502 640574
rect 238586 640338 238822 640574
rect 238266 604658 238502 604894
rect 238586 604658 238822 604894
rect 238266 604338 238502 604574
rect 238586 604338 238822 604574
rect 238266 568658 238502 568894
rect 238586 568658 238822 568894
rect 238266 568338 238502 568574
rect 238586 568338 238822 568574
rect 238266 532658 238502 532894
rect 238586 532658 238822 532894
rect 238266 532338 238502 532574
rect 238586 532338 238822 532574
rect 238266 496658 238502 496894
rect 238586 496658 238822 496894
rect 238266 496338 238502 496574
rect 238586 496338 238822 496574
rect 238266 460658 238502 460894
rect 238586 460658 238822 460894
rect 238266 460338 238502 460574
rect 238586 460338 238822 460574
rect 238266 424658 238502 424894
rect 238586 424658 238822 424894
rect 238266 424338 238502 424574
rect 238586 424338 238822 424574
rect 238266 388658 238502 388894
rect 238586 388658 238822 388894
rect 238266 388338 238502 388574
rect 238586 388338 238822 388574
rect 238266 352658 238502 352894
rect 238586 352658 238822 352894
rect 238266 352338 238502 352574
rect 238586 352338 238822 352574
rect 238266 316658 238502 316894
rect 238586 316658 238822 316894
rect 238266 316338 238502 316574
rect 238586 316338 238822 316574
rect 238266 280658 238502 280894
rect 238586 280658 238822 280894
rect 238266 280338 238502 280574
rect 238586 280338 238822 280574
rect 238266 244658 238502 244894
rect 238586 244658 238822 244894
rect 238266 244338 238502 244574
rect 238586 244338 238822 244574
rect 238266 208658 238502 208894
rect 238586 208658 238822 208894
rect 238266 208338 238502 208574
rect 238586 208338 238822 208574
rect 238266 172658 238502 172894
rect 238586 172658 238822 172894
rect 238266 172338 238502 172574
rect 238586 172338 238822 172574
rect 238266 136658 238502 136894
rect 238586 136658 238822 136894
rect 238266 136338 238502 136574
rect 238586 136338 238822 136574
rect 238266 100658 238502 100894
rect 238586 100658 238822 100894
rect 238266 100338 238502 100574
rect 238586 100338 238822 100574
rect 238266 64658 238502 64894
rect 238586 64658 238822 64894
rect 238266 64338 238502 64574
rect 238586 64338 238822 64574
rect 238266 28658 238502 28894
rect 238586 28658 238822 28894
rect 238266 28338 238502 28574
rect 238586 28338 238822 28574
rect 240826 704602 241062 704838
rect 241146 704602 241382 704838
rect 240826 704282 241062 704518
rect 241146 704282 241382 704518
rect 240826 687218 241062 687454
rect 241146 687218 241382 687454
rect 240826 686898 241062 687134
rect 241146 686898 241382 687134
rect 240826 651218 241062 651454
rect 241146 651218 241382 651454
rect 240826 650898 241062 651134
rect 241146 650898 241382 651134
rect 240826 615218 241062 615454
rect 241146 615218 241382 615454
rect 240826 614898 241062 615134
rect 241146 614898 241382 615134
rect 240826 579218 241062 579454
rect 241146 579218 241382 579454
rect 240826 578898 241062 579134
rect 241146 578898 241382 579134
rect 240826 543218 241062 543454
rect 241146 543218 241382 543454
rect 240826 542898 241062 543134
rect 241146 542898 241382 543134
rect 240826 507218 241062 507454
rect 241146 507218 241382 507454
rect 240826 506898 241062 507134
rect 241146 506898 241382 507134
rect 240826 471218 241062 471454
rect 241146 471218 241382 471454
rect 240826 470898 241062 471134
rect 241146 470898 241382 471134
rect 240826 435218 241062 435454
rect 241146 435218 241382 435454
rect 240826 434898 241062 435134
rect 241146 434898 241382 435134
rect 240826 399218 241062 399454
rect 241146 399218 241382 399454
rect 240826 398898 241062 399134
rect 241146 398898 241382 399134
rect 240826 363218 241062 363454
rect 241146 363218 241382 363454
rect 240826 362898 241062 363134
rect 241146 362898 241382 363134
rect 240826 327218 241062 327454
rect 241146 327218 241382 327454
rect 240826 326898 241062 327134
rect 241146 326898 241382 327134
rect 240826 291218 241062 291454
rect 241146 291218 241382 291454
rect 240826 290898 241062 291134
rect 241146 290898 241382 291134
rect 240826 255218 241062 255454
rect 241146 255218 241382 255454
rect 240826 254898 241062 255134
rect 241146 254898 241382 255134
rect 240826 219218 241062 219454
rect 241146 219218 241382 219454
rect 240826 218898 241062 219134
rect 241146 218898 241382 219134
rect 240826 183218 241062 183454
rect 241146 183218 241382 183454
rect 240826 182898 241062 183134
rect 241146 182898 241382 183134
rect 240826 147218 241062 147454
rect 241146 147218 241382 147454
rect 240826 146898 241062 147134
rect 241146 146898 241382 147134
rect 240826 111218 241062 111454
rect 241146 111218 241382 111454
rect 240826 110898 241062 111134
rect 241146 110898 241382 111134
rect 240826 75218 241062 75454
rect 241146 75218 241382 75454
rect 240826 74898 241062 75134
rect 241146 74898 241382 75134
rect 240826 39218 241062 39454
rect 241146 39218 241382 39454
rect 240826 38898 241062 39134
rect 241146 38898 241382 39134
rect 240826 3218 241062 3454
rect 241146 3218 241382 3454
rect 240826 2898 241062 3134
rect 241146 2898 241382 3134
rect 240826 -582 241062 -346
rect 241146 -582 241382 -346
rect 240826 -902 241062 -666
rect 241146 -902 241382 -666
rect 251986 710362 252222 710598
rect 252306 710362 252542 710598
rect 251986 710042 252222 710278
rect 252306 710042 252542 710278
rect 248266 708442 248502 708678
rect 248586 708442 248822 708678
rect 248266 708122 248502 708358
rect 248586 708122 248822 708358
rect 241986 680378 242222 680614
rect 242306 680378 242542 680614
rect 241986 680058 242222 680294
rect 242306 680058 242542 680294
rect 241986 644378 242222 644614
rect 242306 644378 242542 644614
rect 241986 644058 242222 644294
rect 242306 644058 242542 644294
rect 241986 608378 242222 608614
rect 242306 608378 242542 608614
rect 241986 608058 242222 608294
rect 242306 608058 242542 608294
rect 241986 572378 242222 572614
rect 242306 572378 242542 572614
rect 241986 572058 242222 572294
rect 242306 572058 242542 572294
rect 241986 536378 242222 536614
rect 242306 536378 242542 536614
rect 241986 536058 242222 536294
rect 242306 536058 242542 536294
rect 241986 500378 242222 500614
rect 242306 500378 242542 500614
rect 241986 500058 242222 500294
rect 242306 500058 242542 500294
rect 241986 464378 242222 464614
rect 242306 464378 242542 464614
rect 241986 464058 242222 464294
rect 242306 464058 242542 464294
rect 241986 428378 242222 428614
rect 242306 428378 242542 428614
rect 241986 428058 242222 428294
rect 242306 428058 242542 428294
rect 241986 392378 242222 392614
rect 242306 392378 242542 392614
rect 241986 392058 242222 392294
rect 242306 392058 242542 392294
rect 241986 356378 242222 356614
rect 242306 356378 242542 356614
rect 241986 356058 242222 356294
rect 242306 356058 242542 356294
rect 241986 320378 242222 320614
rect 242306 320378 242542 320614
rect 241986 320058 242222 320294
rect 242306 320058 242542 320294
rect 241986 284378 242222 284614
rect 242306 284378 242542 284614
rect 241986 284058 242222 284294
rect 242306 284058 242542 284294
rect 241986 248378 242222 248614
rect 242306 248378 242542 248614
rect 241986 248058 242222 248294
rect 242306 248058 242542 248294
rect 241986 212378 242222 212614
rect 242306 212378 242542 212614
rect 241986 212058 242222 212294
rect 242306 212058 242542 212294
rect 241986 176378 242222 176614
rect 242306 176378 242542 176614
rect 241986 176058 242222 176294
rect 242306 176058 242542 176294
rect 241986 140378 242222 140614
rect 242306 140378 242542 140614
rect 241986 140058 242222 140294
rect 242306 140058 242542 140294
rect 241986 104378 242222 104614
rect 242306 104378 242542 104614
rect 241986 104058 242222 104294
rect 242306 104058 242542 104294
rect 241986 68378 242222 68614
rect 242306 68378 242542 68614
rect 241986 68058 242222 68294
rect 242306 68058 242542 68294
rect 241986 32378 242222 32614
rect 242306 32378 242542 32614
rect 241986 32058 242222 32294
rect 242306 32058 242542 32294
rect 238266 -5382 238502 -5146
rect 238586 -5382 238822 -5146
rect 238266 -5702 238502 -5466
rect 238586 -5702 238822 -5466
rect 231986 -6342 232222 -6106
rect 232306 -6342 232542 -6106
rect 231986 -6662 232222 -6426
rect 232306 -6662 232542 -6426
rect 244546 706522 244782 706758
rect 244866 706522 245102 706758
rect 244546 706202 244782 706438
rect 244866 706202 245102 706438
rect 244546 690938 244782 691174
rect 244866 690938 245102 691174
rect 244546 690618 244782 690854
rect 244866 690618 245102 690854
rect 244546 654938 244782 655174
rect 244866 654938 245102 655174
rect 244546 654618 244782 654854
rect 244866 654618 245102 654854
rect 244546 618938 244782 619174
rect 244866 618938 245102 619174
rect 244546 618618 244782 618854
rect 244866 618618 245102 618854
rect 244546 582938 244782 583174
rect 244866 582938 245102 583174
rect 244546 582618 244782 582854
rect 244866 582618 245102 582854
rect 244546 546938 244782 547174
rect 244866 546938 245102 547174
rect 244546 546618 244782 546854
rect 244866 546618 245102 546854
rect 244546 510938 244782 511174
rect 244866 510938 245102 511174
rect 244546 510618 244782 510854
rect 244866 510618 245102 510854
rect 244546 474938 244782 475174
rect 244866 474938 245102 475174
rect 244546 474618 244782 474854
rect 244866 474618 245102 474854
rect 244546 438938 244782 439174
rect 244866 438938 245102 439174
rect 244546 438618 244782 438854
rect 244866 438618 245102 438854
rect 244546 402938 244782 403174
rect 244866 402938 245102 403174
rect 244546 402618 244782 402854
rect 244866 402618 245102 402854
rect 244546 366938 244782 367174
rect 244866 366938 245102 367174
rect 244546 366618 244782 366854
rect 244866 366618 245102 366854
rect 244546 330938 244782 331174
rect 244866 330938 245102 331174
rect 244546 330618 244782 330854
rect 244866 330618 245102 330854
rect 244546 294938 244782 295174
rect 244866 294938 245102 295174
rect 244546 294618 244782 294854
rect 244866 294618 245102 294854
rect 244546 258938 244782 259174
rect 244866 258938 245102 259174
rect 244546 258618 244782 258854
rect 244866 258618 245102 258854
rect 244546 222938 244782 223174
rect 244866 222938 245102 223174
rect 244546 222618 244782 222854
rect 244866 222618 245102 222854
rect 244546 186938 244782 187174
rect 244866 186938 245102 187174
rect 244546 186618 244782 186854
rect 244866 186618 245102 186854
rect 244546 150938 244782 151174
rect 244866 150938 245102 151174
rect 244546 150618 244782 150854
rect 244866 150618 245102 150854
rect 244546 114938 244782 115174
rect 244866 114938 245102 115174
rect 244546 114618 244782 114854
rect 244866 114618 245102 114854
rect 244546 78938 244782 79174
rect 244866 78938 245102 79174
rect 244546 78618 244782 78854
rect 244866 78618 245102 78854
rect 244546 42938 244782 43174
rect 244866 42938 245102 43174
rect 244546 42618 244782 42854
rect 244866 42618 245102 42854
rect 244546 6938 244782 7174
rect 244866 6938 245102 7174
rect 244546 6618 244782 6854
rect 244866 6618 245102 6854
rect 244546 -2502 244782 -2266
rect 244866 -2502 245102 -2266
rect 244546 -2822 244782 -2586
rect 244866 -2822 245102 -2586
rect 248266 694658 248502 694894
rect 248586 694658 248822 694894
rect 248266 694338 248502 694574
rect 248586 694338 248822 694574
rect 248266 658658 248502 658894
rect 248586 658658 248822 658894
rect 248266 658338 248502 658574
rect 248586 658338 248822 658574
rect 248266 622658 248502 622894
rect 248586 622658 248822 622894
rect 248266 622338 248502 622574
rect 248586 622338 248822 622574
rect 248266 586658 248502 586894
rect 248586 586658 248822 586894
rect 248266 586338 248502 586574
rect 248586 586338 248822 586574
rect 248266 550658 248502 550894
rect 248586 550658 248822 550894
rect 248266 550338 248502 550574
rect 248586 550338 248822 550574
rect 248266 514658 248502 514894
rect 248586 514658 248822 514894
rect 248266 514338 248502 514574
rect 248586 514338 248822 514574
rect 248266 478658 248502 478894
rect 248586 478658 248822 478894
rect 248266 478338 248502 478574
rect 248586 478338 248822 478574
rect 248266 442658 248502 442894
rect 248586 442658 248822 442894
rect 248266 442338 248502 442574
rect 248586 442338 248822 442574
rect 248266 406658 248502 406894
rect 248586 406658 248822 406894
rect 248266 406338 248502 406574
rect 248586 406338 248822 406574
rect 248266 370658 248502 370894
rect 248586 370658 248822 370894
rect 248266 370338 248502 370574
rect 248586 370338 248822 370574
rect 248266 334658 248502 334894
rect 248586 334658 248822 334894
rect 248266 334338 248502 334574
rect 248586 334338 248822 334574
rect 248266 298658 248502 298894
rect 248586 298658 248822 298894
rect 248266 298338 248502 298574
rect 248586 298338 248822 298574
rect 248266 262658 248502 262894
rect 248586 262658 248822 262894
rect 248266 262338 248502 262574
rect 248586 262338 248822 262574
rect 248266 226658 248502 226894
rect 248586 226658 248822 226894
rect 248266 226338 248502 226574
rect 248586 226338 248822 226574
rect 248266 190658 248502 190894
rect 248586 190658 248822 190894
rect 248266 190338 248502 190574
rect 248586 190338 248822 190574
rect 248266 154658 248502 154894
rect 248586 154658 248822 154894
rect 248266 154338 248502 154574
rect 248586 154338 248822 154574
rect 248266 118658 248502 118894
rect 248586 118658 248822 118894
rect 248266 118338 248502 118574
rect 248586 118338 248822 118574
rect 248266 82658 248502 82894
rect 248586 82658 248822 82894
rect 248266 82338 248502 82574
rect 248586 82338 248822 82574
rect 248266 46658 248502 46894
rect 248586 46658 248822 46894
rect 248266 46338 248502 46574
rect 248586 46338 248822 46574
rect 248266 10658 248502 10894
rect 248586 10658 248822 10894
rect 248266 10338 248502 10574
rect 248586 10338 248822 10574
rect 250826 705562 251062 705798
rect 251146 705562 251382 705798
rect 250826 705242 251062 705478
rect 251146 705242 251382 705478
rect 250826 669218 251062 669454
rect 251146 669218 251382 669454
rect 250826 668898 251062 669134
rect 251146 668898 251382 669134
rect 250826 633218 251062 633454
rect 251146 633218 251382 633454
rect 250826 632898 251062 633134
rect 251146 632898 251382 633134
rect 250826 597218 251062 597454
rect 251146 597218 251382 597454
rect 250826 596898 251062 597134
rect 251146 596898 251382 597134
rect 250826 561218 251062 561454
rect 251146 561218 251382 561454
rect 250826 560898 251062 561134
rect 251146 560898 251382 561134
rect 250826 525218 251062 525454
rect 251146 525218 251382 525454
rect 250826 524898 251062 525134
rect 251146 524898 251382 525134
rect 250826 489218 251062 489454
rect 251146 489218 251382 489454
rect 250826 488898 251062 489134
rect 251146 488898 251382 489134
rect 250826 453218 251062 453454
rect 251146 453218 251382 453454
rect 250826 452898 251062 453134
rect 251146 452898 251382 453134
rect 250826 417218 251062 417454
rect 251146 417218 251382 417454
rect 250826 416898 251062 417134
rect 251146 416898 251382 417134
rect 250826 381218 251062 381454
rect 251146 381218 251382 381454
rect 250826 380898 251062 381134
rect 251146 380898 251382 381134
rect 250826 345218 251062 345454
rect 251146 345218 251382 345454
rect 250826 344898 251062 345134
rect 251146 344898 251382 345134
rect 250826 309218 251062 309454
rect 251146 309218 251382 309454
rect 250826 308898 251062 309134
rect 251146 308898 251382 309134
rect 250826 273218 251062 273454
rect 251146 273218 251382 273454
rect 250826 272898 251062 273134
rect 251146 272898 251382 273134
rect 250826 237218 251062 237454
rect 251146 237218 251382 237454
rect 250826 236898 251062 237134
rect 251146 236898 251382 237134
rect 250826 201218 251062 201454
rect 251146 201218 251382 201454
rect 250826 200898 251062 201134
rect 251146 200898 251382 201134
rect 250826 165218 251062 165454
rect 251146 165218 251382 165454
rect 250826 164898 251062 165134
rect 251146 164898 251382 165134
rect 250826 129218 251062 129454
rect 251146 129218 251382 129454
rect 250826 128898 251062 129134
rect 251146 128898 251382 129134
rect 250826 93218 251062 93454
rect 251146 93218 251382 93454
rect 250826 92898 251062 93134
rect 251146 92898 251382 93134
rect 250826 57218 251062 57454
rect 251146 57218 251382 57454
rect 250826 56898 251062 57134
rect 251146 56898 251382 57134
rect 250826 21218 251062 21454
rect 251146 21218 251382 21454
rect 250826 20898 251062 21134
rect 251146 20898 251382 21134
rect 250826 -1542 251062 -1306
rect 251146 -1542 251382 -1306
rect 250826 -1862 251062 -1626
rect 251146 -1862 251382 -1626
rect 261986 711322 262222 711558
rect 262306 711322 262542 711558
rect 261986 711002 262222 711238
rect 262306 711002 262542 711238
rect 258266 709402 258502 709638
rect 258586 709402 258822 709638
rect 258266 709082 258502 709318
rect 258586 709082 258822 709318
rect 251986 698378 252222 698614
rect 252306 698378 252542 698614
rect 251986 698058 252222 698294
rect 252306 698058 252542 698294
rect 251986 662378 252222 662614
rect 252306 662378 252542 662614
rect 251986 662058 252222 662294
rect 252306 662058 252542 662294
rect 251986 626378 252222 626614
rect 252306 626378 252542 626614
rect 251986 626058 252222 626294
rect 252306 626058 252542 626294
rect 251986 590378 252222 590614
rect 252306 590378 252542 590614
rect 251986 590058 252222 590294
rect 252306 590058 252542 590294
rect 251986 554378 252222 554614
rect 252306 554378 252542 554614
rect 251986 554058 252222 554294
rect 252306 554058 252542 554294
rect 251986 518378 252222 518614
rect 252306 518378 252542 518614
rect 251986 518058 252222 518294
rect 252306 518058 252542 518294
rect 251986 482378 252222 482614
rect 252306 482378 252542 482614
rect 251986 482058 252222 482294
rect 252306 482058 252542 482294
rect 251986 446378 252222 446614
rect 252306 446378 252542 446614
rect 251986 446058 252222 446294
rect 252306 446058 252542 446294
rect 251986 410378 252222 410614
rect 252306 410378 252542 410614
rect 251986 410058 252222 410294
rect 252306 410058 252542 410294
rect 251986 374378 252222 374614
rect 252306 374378 252542 374614
rect 251986 374058 252222 374294
rect 252306 374058 252542 374294
rect 251986 338378 252222 338614
rect 252306 338378 252542 338614
rect 251986 338058 252222 338294
rect 252306 338058 252542 338294
rect 251986 302378 252222 302614
rect 252306 302378 252542 302614
rect 251986 302058 252222 302294
rect 252306 302058 252542 302294
rect 251986 266378 252222 266614
rect 252306 266378 252542 266614
rect 251986 266058 252222 266294
rect 252306 266058 252542 266294
rect 251986 230378 252222 230614
rect 252306 230378 252542 230614
rect 251986 230058 252222 230294
rect 252306 230058 252542 230294
rect 251986 194378 252222 194614
rect 252306 194378 252542 194614
rect 251986 194058 252222 194294
rect 252306 194058 252542 194294
rect 251986 158378 252222 158614
rect 252306 158378 252542 158614
rect 251986 158058 252222 158294
rect 252306 158058 252542 158294
rect 251986 122378 252222 122614
rect 252306 122378 252542 122614
rect 251986 122058 252222 122294
rect 252306 122058 252542 122294
rect 251986 86378 252222 86614
rect 252306 86378 252542 86614
rect 251986 86058 252222 86294
rect 252306 86058 252542 86294
rect 251986 50378 252222 50614
rect 252306 50378 252542 50614
rect 251986 50058 252222 50294
rect 252306 50058 252542 50294
rect 251986 14378 252222 14614
rect 252306 14378 252542 14614
rect 251986 14058 252222 14294
rect 252306 14058 252542 14294
rect 248266 -4422 248502 -4186
rect 248586 -4422 248822 -4186
rect 248266 -4742 248502 -4506
rect 248586 -4742 248822 -4506
rect 241986 -7302 242222 -7066
rect 242306 -7302 242542 -7066
rect 241986 -7622 242222 -7386
rect 242306 -7622 242542 -7386
rect 254546 707482 254782 707718
rect 254866 707482 255102 707718
rect 254546 707162 254782 707398
rect 254866 707162 255102 707398
rect 254546 672938 254782 673174
rect 254866 672938 255102 673174
rect 254546 672618 254782 672854
rect 254866 672618 255102 672854
rect 254546 636938 254782 637174
rect 254866 636938 255102 637174
rect 254546 636618 254782 636854
rect 254866 636618 255102 636854
rect 254546 600938 254782 601174
rect 254866 600938 255102 601174
rect 254546 600618 254782 600854
rect 254866 600618 255102 600854
rect 254546 564938 254782 565174
rect 254866 564938 255102 565174
rect 254546 564618 254782 564854
rect 254866 564618 255102 564854
rect 254546 528938 254782 529174
rect 254866 528938 255102 529174
rect 254546 528618 254782 528854
rect 254866 528618 255102 528854
rect 254546 492938 254782 493174
rect 254866 492938 255102 493174
rect 254546 492618 254782 492854
rect 254866 492618 255102 492854
rect 254546 456938 254782 457174
rect 254866 456938 255102 457174
rect 254546 456618 254782 456854
rect 254866 456618 255102 456854
rect 254546 420938 254782 421174
rect 254866 420938 255102 421174
rect 254546 420618 254782 420854
rect 254866 420618 255102 420854
rect 254546 384938 254782 385174
rect 254866 384938 255102 385174
rect 254546 384618 254782 384854
rect 254866 384618 255102 384854
rect 254546 348938 254782 349174
rect 254866 348938 255102 349174
rect 254546 348618 254782 348854
rect 254866 348618 255102 348854
rect 254546 312938 254782 313174
rect 254866 312938 255102 313174
rect 254546 312618 254782 312854
rect 254866 312618 255102 312854
rect 254546 276938 254782 277174
rect 254866 276938 255102 277174
rect 254546 276618 254782 276854
rect 254866 276618 255102 276854
rect 254546 240938 254782 241174
rect 254866 240938 255102 241174
rect 254546 240618 254782 240854
rect 254866 240618 255102 240854
rect 254546 204938 254782 205174
rect 254866 204938 255102 205174
rect 254546 204618 254782 204854
rect 254866 204618 255102 204854
rect 254546 168938 254782 169174
rect 254866 168938 255102 169174
rect 254546 168618 254782 168854
rect 254866 168618 255102 168854
rect 254546 132938 254782 133174
rect 254866 132938 255102 133174
rect 254546 132618 254782 132854
rect 254866 132618 255102 132854
rect 254546 96938 254782 97174
rect 254866 96938 255102 97174
rect 254546 96618 254782 96854
rect 254866 96618 255102 96854
rect 254546 60938 254782 61174
rect 254866 60938 255102 61174
rect 254546 60618 254782 60854
rect 254866 60618 255102 60854
rect 254546 24938 254782 25174
rect 254866 24938 255102 25174
rect 254546 24618 254782 24854
rect 254866 24618 255102 24854
rect 254546 -3462 254782 -3226
rect 254866 -3462 255102 -3226
rect 254546 -3782 254782 -3546
rect 254866 -3782 255102 -3546
rect 258266 676658 258502 676894
rect 258586 676658 258822 676894
rect 258266 676338 258502 676574
rect 258586 676338 258822 676574
rect 258266 640658 258502 640894
rect 258586 640658 258822 640894
rect 258266 640338 258502 640574
rect 258586 640338 258822 640574
rect 258266 604658 258502 604894
rect 258586 604658 258822 604894
rect 258266 604338 258502 604574
rect 258586 604338 258822 604574
rect 258266 568658 258502 568894
rect 258586 568658 258822 568894
rect 258266 568338 258502 568574
rect 258586 568338 258822 568574
rect 258266 532658 258502 532894
rect 258586 532658 258822 532894
rect 258266 532338 258502 532574
rect 258586 532338 258822 532574
rect 258266 496658 258502 496894
rect 258586 496658 258822 496894
rect 258266 496338 258502 496574
rect 258586 496338 258822 496574
rect 258266 460658 258502 460894
rect 258586 460658 258822 460894
rect 258266 460338 258502 460574
rect 258586 460338 258822 460574
rect 258266 424658 258502 424894
rect 258586 424658 258822 424894
rect 258266 424338 258502 424574
rect 258586 424338 258822 424574
rect 258266 388658 258502 388894
rect 258586 388658 258822 388894
rect 258266 388338 258502 388574
rect 258586 388338 258822 388574
rect 258266 352658 258502 352894
rect 258586 352658 258822 352894
rect 258266 352338 258502 352574
rect 258586 352338 258822 352574
rect 258266 316658 258502 316894
rect 258586 316658 258822 316894
rect 258266 316338 258502 316574
rect 258586 316338 258822 316574
rect 258266 280658 258502 280894
rect 258586 280658 258822 280894
rect 258266 280338 258502 280574
rect 258586 280338 258822 280574
rect 258266 244658 258502 244894
rect 258586 244658 258822 244894
rect 258266 244338 258502 244574
rect 258586 244338 258822 244574
rect 258266 208658 258502 208894
rect 258586 208658 258822 208894
rect 258266 208338 258502 208574
rect 258586 208338 258822 208574
rect 258266 172658 258502 172894
rect 258586 172658 258822 172894
rect 258266 172338 258502 172574
rect 258586 172338 258822 172574
rect 258266 136658 258502 136894
rect 258586 136658 258822 136894
rect 258266 136338 258502 136574
rect 258586 136338 258822 136574
rect 258266 100658 258502 100894
rect 258586 100658 258822 100894
rect 258266 100338 258502 100574
rect 258586 100338 258822 100574
rect 258266 64658 258502 64894
rect 258586 64658 258822 64894
rect 258266 64338 258502 64574
rect 258586 64338 258822 64574
rect 258266 28658 258502 28894
rect 258586 28658 258822 28894
rect 258266 28338 258502 28574
rect 258586 28338 258822 28574
rect 260826 704602 261062 704838
rect 261146 704602 261382 704838
rect 260826 704282 261062 704518
rect 261146 704282 261382 704518
rect 260826 687218 261062 687454
rect 261146 687218 261382 687454
rect 260826 686898 261062 687134
rect 261146 686898 261382 687134
rect 260826 651218 261062 651454
rect 261146 651218 261382 651454
rect 260826 650898 261062 651134
rect 261146 650898 261382 651134
rect 260826 615218 261062 615454
rect 261146 615218 261382 615454
rect 260826 614898 261062 615134
rect 261146 614898 261382 615134
rect 260826 579218 261062 579454
rect 261146 579218 261382 579454
rect 260826 578898 261062 579134
rect 261146 578898 261382 579134
rect 260826 543218 261062 543454
rect 261146 543218 261382 543454
rect 260826 542898 261062 543134
rect 261146 542898 261382 543134
rect 260826 507218 261062 507454
rect 261146 507218 261382 507454
rect 260826 506898 261062 507134
rect 261146 506898 261382 507134
rect 260826 471218 261062 471454
rect 261146 471218 261382 471454
rect 260826 470898 261062 471134
rect 261146 470898 261382 471134
rect 260826 435218 261062 435454
rect 261146 435218 261382 435454
rect 260826 434898 261062 435134
rect 261146 434898 261382 435134
rect 260826 399218 261062 399454
rect 261146 399218 261382 399454
rect 260826 398898 261062 399134
rect 261146 398898 261382 399134
rect 260826 363218 261062 363454
rect 261146 363218 261382 363454
rect 260826 362898 261062 363134
rect 261146 362898 261382 363134
rect 260826 327218 261062 327454
rect 261146 327218 261382 327454
rect 260826 326898 261062 327134
rect 261146 326898 261382 327134
rect 260826 291218 261062 291454
rect 261146 291218 261382 291454
rect 260826 290898 261062 291134
rect 261146 290898 261382 291134
rect 260826 255218 261062 255454
rect 261146 255218 261382 255454
rect 260826 254898 261062 255134
rect 261146 254898 261382 255134
rect 260826 219218 261062 219454
rect 261146 219218 261382 219454
rect 260826 218898 261062 219134
rect 261146 218898 261382 219134
rect 260826 183218 261062 183454
rect 261146 183218 261382 183454
rect 260826 182898 261062 183134
rect 261146 182898 261382 183134
rect 260826 147218 261062 147454
rect 261146 147218 261382 147454
rect 260826 146898 261062 147134
rect 261146 146898 261382 147134
rect 260826 111218 261062 111454
rect 261146 111218 261382 111454
rect 260826 110898 261062 111134
rect 261146 110898 261382 111134
rect 260826 75218 261062 75454
rect 261146 75218 261382 75454
rect 260826 74898 261062 75134
rect 261146 74898 261382 75134
rect 260826 39218 261062 39454
rect 261146 39218 261382 39454
rect 260826 38898 261062 39134
rect 261146 38898 261382 39134
rect 260826 3218 261062 3454
rect 261146 3218 261382 3454
rect 260826 2898 261062 3134
rect 261146 2898 261382 3134
rect 260826 -582 261062 -346
rect 261146 -582 261382 -346
rect 260826 -902 261062 -666
rect 261146 -902 261382 -666
rect 271986 710362 272222 710598
rect 272306 710362 272542 710598
rect 271986 710042 272222 710278
rect 272306 710042 272542 710278
rect 268266 708442 268502 708678
rect 268586 708442 268822 708678
rect 268266 708122 268502 708358
rect 268586 708122 268822 708358
rect 261986 680378 262222 680614
rect 262306 680378 262542 680614
rect 261986 680058 262222 680294
rect 262306 680058 262542 680294
rect 261986 644378 262222 644614
rect 262306 644378 262542 644614
rect 261986 644058 262222 644294
rect 262306 644058 262542 644294
rect 261986 608378 262222 608614
rect 262306 608378 262542 608614
rect 261986 608058 262222 608294
rect 262306 608058 262542 608294
rect 261986 572378 262222 572614
rect 262306 572378 262542 572614
rect 261986 572058 262222 572294
rect 262306 572058 262542 572294
rect 261986 536378 262222 536614
rect 262306 536378 262542 536614
rect 261986 536058 262222 536294
rect 262306 536058 262542 536294
rect 261986 500378 262222 500614
rect 262306 500378 262542 500614
rect 261986 500058 262222 500294
rect 262306 500058 262542 500294
rect 261986 464378 262222 464614
rect 262306 464378 262542 464614
rect 261986 464058 262222 464294
rect 262306 464058 262542 464294
rect 261986 428378 262222 428614
rect 262306 428378 262542 428614
rect 261986 428058 262222 428294
rect 262306 428058 262542 428294
rect 261986 392378 262222 392614
rect 262306 392378 262542 392614
rect 261986 392058 262222 392294
rect 262306 392058 262542 392294
rect 261986 356378 262222 356614
rect 262306 356378 262542 356614
rect 261986 356058 262222 356294
rect 262306 356058 262542 356294
rect 261986 320378 262222 320614
rect 262306 320378 262542 320614
rect 261986 320058 262222 320294
rect 262306 320058 262542 320294
rect 261986 284378 262222 284614
rect 262306 284378 262542 284614
rect 261986 284058 262222 284294
rect 262306 284058 262542 284294
rect 261986 248378 262222 248614
rect 262306 248378 262542 248614
rect 261986 248058 262222 248294
rect 262306 248058 262542 248294
rect 261986 212378 262222 212614
rect 262306 212378 262542 212614
rect 261986 212058 262222 212294
rect 262306 212058 262542 212294
rect 261986 176378 262222 176614
rect 262306 176378 262542 176614
rect 261986 176058 262222 176294
rect 262306 176058 262542 176294
rect 261986 140378 262222 140614
rect 262306 140378 262542 140614
rect 261986 140058 262222 140294
rect 262306 140058 262542 140294
rect 261986 104378 262222 104614
rect 262306 104378 262542 104614
rect 261986 104058 262222 104294
rect 262306 104058 262542 104294
rect 261986 68378 262222 68614
rect 262306 68378 262542 68614
rect 261986 68058 262222 68294
rect 262306 68058 262542 68294
rect 261986 32378 262222 32614
rect 262306 32378 262542 32614
rect 261986 32058 262222 32294
rect 262306 32058 262542 32294
rect 258266 -5382 258502 -5146
rect 258586 -5382 258822 -5146
rect 258266 -5702 258502 -5466
rect 258586 -5702 258822 -5466
rect 251986 -6342 252222 -6106
rect 252306 -6342 252542 -6106
rect 251986 -6662 252222 -6426
rect 252306 -6662 252542 -6426
rect 264546 706522 264782 706758
rect 264866 706522 265102 706758
rect 264546 706202 264782 706438
rect 264866 706202 265102 706438
rect 264546 690938 264782 691174
rect 264866 690938 265102 691174
rect 264546 690618 264782 690854
rect 264866 690618 265102 690854
rect 264546 654938 264782 655174
rect 264866 654938 265102 655174
rect 264546 654618 264782 654854
rect 264866 654618 265102 654854
rect 264546 618938 264782 619174
rect 264866 618938 265102 619174
rect 264546 618618 264782 618854
rect 264866 618618 265102 618854
rect 264546 582938 264782 583174
rect 264866 582938 265102 583174
rect 264546 582618 264782 582854
rect 264866 582618 265102 582854
rect 264546 546938 264782 547174
rect 264866 546938 265102 547174
rect 264546 546618 264782 546854
rect 264866 546618 265102 546854
rect 264546 510938 264782 511174
rect 264866 510938 265102 511174
rect 264546 510618 264782 510854
rect 264866 510618 265102 510854
rect 264546 474938 264782 475174
rect 264866 474938 265102 475174
rect 264546 474618 264782 474854
rect 264866 474618 265102 474854
rect 264546 438938 264782 439174
rect 264866 438938 265102 439174
rect 264546 438618 264782 438854
rect 264866 438618 265102 438854
rect 264546 402938 264782 403174
rect 264866 402938 265102 403174
rect 264546 402618 264782 402854
rect 264866 402618 265102 402854
rect 264546 366938 264782 367174
rect 264866 366938 265102 367174
rect 264546 366618 264782 366854
rect 264866 366618 265102 366854
rect 264546 330938 264782 331174
rect 264866 330938 265102 331174
rect 264546 330618 264782 330854
rect 264866 330618 265102 330854
rect 264546 294938 264782 295174
rect 264866 294938 265102 295174
rect 264546 294618 264782 294854
rect 264866 294618 265102 294854
rect 264546 258938 264782 259174
rect 264866 258938 265102 259174
rect 264546 258618 264782 258854
rect 264866 258618 265102 258854
rect 264546 222938 264782 223174
rect 264866 222938 265102 223174
rect 264546 222618 264782 222854
rect 264866 222618 265102 222854
rect 264546 186938 264782 187174
rect 264866 186938 265102 187174
rect 264546 186618 264782 186854
rect 264866 186618 265102 186854
rect 264546 150938 264782 151174
rect 264866 150938 265102 151174
rect 264546 150618 264782 150854
rect 264866 150618 265102 150854
rect 264546 114938 264782 115174
rect 264866 114938 265102 115174
rect 264546 114618 264782 114854
rect 264866 114618 265102 114854
rect 264546 78938 264782 79174
rect 264866 78938 265102 79174
rect 264546 78618 264782 78854
rect 264866 78618 265102 78854
rect 264546 42938 264782 43174
rect 264866 42938 265102 43174
rect 264546 42618 264782 42854
rect 264866 42618 265102 42854
rect 264546 6938 264782 7174
rect 264866 6938 265102 7174
rect 264546 6618 264782 6854
rect 264866 6618 265102 6854
rect 264546 -2502 264782 -2266
rect 264866 -2502 265102 -2266
rect 264546 -2822 264782 -2586
rect 264866 -2822 265102 -2586
rect 268266 694658 268502 694894
rect 268586 694658 268822 694894
rect 268266 694338 268502 694574
rect 268586 694338 268822 694574
rect 268266 658658 268502 658894
rect 268586 658658 268822 658894
rect 268266 658338 268502 658574
rect 268586 658338 268822 658574
rect 268266 622658 268502 622894
rect 268586 622658 268822 622894
rect 268266 622338 268502 622574
rect 268586 622338 268822 622574
rect 268266 586658 268502 586894
rect 268586 586658 268822 586894
rect 268266 586338 268502 586574
rect 268586 586338 268822 586574
rect 268266 550658 268502 550894
rect 268586 550658 268822 550894
rect 268266 550338 268502 550574
rect 268586 550338 268822 550574
rect 268266 514658 268502 514894
rect 268586 514658 268822 514894
rect 268266 514338 268502 514574
rect 268586 514338 268822 514574
rect 268266 478658 268502 478894
rect 268586 478658 268822 478894
rect 268266 478338 268502 478574
rect 268586 478338 268822 478574
rect 268266 442658 268502 442894
rect 268586 442658 268822 442894
rect 268266 442338 268502 442574
rect 268586 442338 268822 442574
rect 268266 406658 268502 406894
rect 268586 406658 268822 406894
rect 268266 406338 268502 406574
rect 268586 406338 268822 406574
rect 268266 370658 268502 370894
rect 268586 370658 268822 370894
rect 268266 370338 268502 370574
rect 268586 370338 268822 370574
rect 268266 334658 268502 334894
rect 268586 334658 268822 334894
rect 268266 334338 268502 334574
rect 268586 334338 268822 334574
rect 268266 298658 268502 298894
rect 268586 298658 268822 298894
rect 268266 298338 268502 298574
rect 268586 298338 268822 298574
rect 268266 262658 268502 262894
rect 268586 262658 268822 262894
rect 268266 262338 268502 262574
rect 268586 262338 268822 262574
rect 268266 226658 268502 226894
rect 268586 226658 268822 226894
rect 268266 226338 268502 226574
rect 268586 226338 268822 226574
rect 268266 190658 268502 190894
rect 268586 190658 268822 190894
rect 268266 190338 268502 190574
rect 268586 190338 268822 190574
rect 268266 154658 268502 154894
rect 268586 154658 268822 154894
rect 268266 154338 268502 154574
rect 268586 154338 268822 154574
rect 268266 118658 268502 118894
rect 268586 118658 268822 118894
rect 268266 118338 268502 118574
rect 268586 118338 268822 118574
rect 268266 82658 268502 82894
rect 268586 82658 268822 82894
rect 268266 82338 268502 82574
rect 268586 82338 268822 82574
rect 268266 46658 268502 46894
rect 268586 46658 268822 46894
rect 268266 46338 268502 46574
rect 268586 46338 268822 46574
rect 268266 10658 268502 10894
rect 268586 10658 268822 10894
rect 268266 10338 268502 10574
rect 268586 10338 268822 10574
rect 270826 705562 271062 705798
rect 271146 705562 271382 705798
rect 270826 705242 271062 705478
rect 271146 705242 271382 705478
rect 270826 669218 271062 669454
rect 271146 669218 271382 669454
rect 270826 668898 271062 669134
rect 271146 668898 271382 669134
rect 270826 633218 271062 633454
rect 271146 633218 271382 633454
rect 270826 632898 271062 633134
rect 271146 632898 271382 633134
rect 270826 597218 271062 597454
rect 271146 597218 271382 597454
rect 270826 596898 271062 597134
rect 271146 596898 271382 597134
rect 270826 561218 271062 561454
rect 271146 561218 271382 561454
rect 270826 560898 271062 561134
rect 271146 560898 271382 561134
rect 270826 525218 271062 525454
rect 271146 525218 271382 525454
rect 270826 524898 271062 525134
rect 271146 524898 271382 525134
rect 270826 489218 271062 489454
rect 271146 489218 271382 489454
rect 270826 488898 271062 489134
rect 271146 488898 271382 489134
rect 270826 453218 271062 453454
rect 271146 453218 271382 453454
rect 270826 452898 271062 453134
rect 271146 452898 271382 453134
rect 270826 417218 271062 417454
rect 271146 417218 271382 417454
rect 270826 416898 271062 417134
rect 271146 416898 271382 417134
rect 270826 381218 271062 381454
rect 271146 381218 271382 381454
rect 270826 380898 271062 381134
rect 271146 380898 271382 381134
rect 270826 345218 271062 345454
rect 271146 345218 271382 345454
rect 270826 344898 271062 345134
rect 271146 344898 271382 345134
rect 270826 309218 271062 309454
rect 271146 309218 271382 309454
rect 270826 308898 271062 309134
rect 271146 308898 271382 309134
rect 270826 273218 271062 273454
rect 271146 273218 271382 273454
rect 270826 272898 271062 273134
rect 271146 272898 271382 273134
rect 270826 237218 271062 237454
rect 271146 237218 271382 237454
rect 270826 236898 271062 237134
rect 271146 236898 271382 237134
rect 270826 201218 271062 201454
rect 271146 201218 271382 201454
rect 270826 200898 271062 201134
rect 271146 200898 271382 201134
rect 270826 165218 271062 165454
rect 271146 165218 271382 165454
rect 270826 164898 271062 165134
rect 271146 164898 271382 165134
rect 270826 129218 271062 129454
rect 271146 129218 271382 129454
rect 270826 128898 271062 129134
rect 271146 128898 271382 129134
rect 270826 93218 271062 93454
rect 271146 93218 271382 93454
rect 270826 92898 271062 93134
rect 271146 92898 271382 93134
rect 270826 57218 271062 57454
rect 271146 57218 271382 57454
rect 270826 56898 271062 57134
rect 271146 56898 271382 57134
rect 270826 21218 271062 21454
rect 271146 21218 271382 21454
rect 270826 20898 271062 21134
rect 271146 20898 271382 21134
rect 270826 -1542 271062 -1306
rect 271146 -1542 271382 -1306
rect 270826 -1862 271062 -1626
rect 271146 -1862 271382 -1626
rect 281986 711322 282222 711558
rect 282306 711322 282542 711558
rect 281986 711002 282222 711238
rect 282306 711002 282542 711238
rect 278266 709402 278502 709638
rect 278586 709402 278822 709638
rect 278266 709082 278502 709318
rect 278586 709082 278822 709318
rect 271986 698378 272222 698614
rect 272306 698378 272542 698614
rect 271986 698058 272222 698294
rect 272306 698058 272542 698294
rect 271986 662378 272222 662614
rect 272306 662378 272542 662614
rect 271986 662058 272222 662294
rect 272306 662058 272542 662294
rect 271986 626378 272222 626614
rect 272306 626378 272542 626614
rect 271986 626058 272222 626294
rect 272306 626058 272542 626294
rect 271986 590378 272222 590614
rect 272306 590378 272542 590614
rect 271986 590058 272222 590294
rect 272306 590058 272542 590294
rect 271986 554378 272222 554614
rect 272306 554378 272542 554614
rect 271986 554058 272222 554294
rect 272306 554058 272542 554294
rect 271986 518378 272222 518614
rect 272306 518378 272542 518614
rect 271986 518058 272222 518294
rect 272306 518058 272542 518294
rect 271986 482378 272222 482614
rect 272306 482378 272542 482614
rect 271986 482058 272222 482294
rect 272306 482058 272542 482294
rect 271986 446378 272222 446614
rect 272306 446378 272542 446614
rect 271986 446058 272222 446294
rect 272306 446058 272542 446294
rect 271986 410378 272222 410614
rect 272306 410378 272542 410614
rect 271986 410058 272222 410294
rect 272306 410058 272542 410294
rect 271986 374378 272222 374614
rect 272306 374378 272542 374614
rect 271986 374058 272222 374294
rect 272306 374058 272542 374294
rect 271986 338378 272222 338614
rect 272306 338378 272542 338614
rect 271986 338058 272222 338294
rect 272306 338058 272542 338294
rect 271986 302378 272222 302614
rect 272306 302378 272542 302614
rect 271986 302058 272222 302294
rect 272306 302058 272542 302294
rect 271986 266378 272222 266614
rect 272306 266378 272542 266614
rect 271986 266058 272222 266294
rect 272306 266058 272542 266294
rect 271986 230378 272222 230614
rect 272306 230378 272542 230614
rect 271986 230058 272222 230294
rect 272306 230058 272542 230294
rect 271986 194378 272222 194614
rect 272306 194378 272542 194614
rect 271986 194058 272222 194294
rect 272306 194058 272542 194294
rect 271986 158378 272222 158614
rect 272306 158378 272542 158614
rect 271986 158058 272222 158294
rect 272306 158058 272542 158294
rect 271986 122378 272222 122614
rect 272306 122378 272542 122614
rect 271986 122058 272222 122294
rect 272306 122058 272542 122294
rect 271986 86378 272222 86614
rect 272306 86378 272542 86614
rect 271986 86058 272222 86294
rect 272306 86058 272542 86294
rect 271986 50378 272222 50614
rect 272306 50378 272542 50614
rect 271986 50058 272222 50294
rect 272306 50058 272542 50294
rect 271986 14378 272222 14614
rect 272306 14378 272542 14614
rect 271986 14058 272222 14294
rect 272306 14058 272542 14294
rect 268266 -4422 268502 -4186
rect 268586 -4422 268822 -4186
rect 268266 -4742 268502 -4506
rect 268586 -4742 268822 -4506
rect 261986 -7302 262222 -7066
rect 262306 -7302 262542 -7066
rect 261986 -7622 262222 -7386
rect 262306 -7622 262542 -7386
rect 274546 707482 274782 707718
rect 274866 707482 275102 707718
rect 274546 707162 274782 707398
rect 274866 707162 275102 707398
rect 274546 672938 274782 673174
rect 274866 672938 275102 673174
rect 274546 672618 274782 672854
rect 274866 672618 275102 672854
rect 274546 636938 274782 637174
rect 274866 636938 275102 637174
rect 274546 636618 274782 636854
rect 274866 636618 275102 636854
rect 274546 600938 274782 601174
rect 274866 600938 275102 601174
rect 274546 600618 274782 600854
rect 274866 600618 275102 600854
rect 274546 564938 274782 565174
rect 274866 564938 275102 565174
rect 274546 564618 274782 564854
rect 274866 564618 275102 564854
rect 274546 528938 274782 529174
rect 274866 528938 275102 529174
rect 274546 528618 274782 528854
rect 274866 528618 275102 528854
rect 274546 492938 274782 493174
rect 274866 492938 275102 493174
rect 274546 492618 274782 492854
rect 274866 492618 275102 492854
rect 274546 456938 274782 457174
rect 274866 456938 275102 457174
rect 274546 456618 274782 456854
rect 274866 456618 275102 456854
rect 274546 420938 274782 421174
rect 274866 420938 275102 421174
rect 274546 420618 274782 420854
rect 274866 420618 275102 420854
rect 274546 384938 274782 385174
rect 274866 384938 275102 385174
rect 274546 384618 274782 384854
rect 274866 384618 275102 384854
rect 274546 348938 274782 349174
rect 274866 348938 275102 349174
rect 274546 348618 274782 348854
rect 274866 348618 275102 348854
rect 274546 312938 274782 313174
rect 274866 312938 275102 313174
rect 274546 312618 274782 312854
rect 274866 312618 275102 312854
rect 274546 276938 274782 277174
rect 274866 276938 275102 277174
rect 274546 276618 274782 276854
rect 274866 276618 275102 276854
rect 274546 240938 274782 241174
rect 274866 240938 275102 241174
rect 274546 240618 274782 240854
rect 274866 240618 275102 240854
rect 274546 204938 274782 205174
rect 274866 204938 275102 205174
rect 274546 204618 274782 204854
rect 274866 204618 275102 204854
rect 274546 168938 274782 169174
rect 274866 168938 275102 169174
rect 274546 168618 274782 168854
rect 274866 168618 275102 168854
rect 274546 132938 274782 133174
rect 274866 132938 275102 133174
rect 274546 132618 274782 132854
rect 274866 132618 275102 132854
rect 274546 96938 274782 97174
rect 274866 96938 275102 97174
rect 274546 96618 274782 96854
rect 274866 96618 275102 96854
rect 274546 60938 274782 61174
rect 274866 60938 275102 61174
rect 274546 60618 274782 60854
rect 274866 60618 275102 60854
rect 274546 24938 274782 25174
rect 274866 24938 275102 25174
rect 274546 24618 274782 24854
rect 274866 24618 275102 24854
rect 274546 -3462 274782 -3226
rect 274866 -3462 275102 -3226
rect 274546 -3782 274782 -3546
rect 274866 -3782 275102 -3546
rect 278266 676658 278502 676894
rect 278586 676658 278822 676894
rect 278266 676338 278502 676574
rect 278586 676338 278822 676574
rect 278266 640658 278502 640894
rect 278586 640658 278822 640894
rect 278266 640338 278502 640574
rect 278586 640338 278822 640574
rect 278266 604658 278502 604894
rect 278586 604658 278822 604894
rect 278266 604338 278502 604574
rect 278586 604338 278822 604574
rect 278266 568658 278502 568894
rect 278586 568658 278822 568894
rect 278266 568338 278502 568574
rect 278586 568338 278822 568574
rect 278266 532658 278502 532894
rect 278586 532658 278822 532894
rect 278266 532338 278502 532574
rect 278586 532338 278822 532574
rect 278266 496658 278502 496894
rect 278586 496658 278822 496894
rect 278266 496338 278502 496574
rect 278586 496338 278822 496574
rect 278266 460658 278502 460894
rect 278586 460658 278822 460894
rect 278266 460338 278502 460574
rect 278586 460338 278822 460574
rect 278266 424658 278502 424894
rect 278586 424658 278822 424894
rect 278266 424338 278502 424574
rect 278586 424338 278822 424574
rect 278266 388658 278502 388894
rect 278586 388658 278822 388894
rect 278266 388338 278502 388574
rect 278586 388338 278822 388574
rect 278266 352658 278502 352894
rect 278586 352658 278822 352894
rect 278266 352338 278502 352574
rect 278586 352338 278822 352574
rect 278266 316658 278502 316894
rect 278586 316658 278822 316894
rect 278266 316338 278502 316574
rect 278586 316338 278822 316574
rect 278266 280658 278502 280894
rect 278586 280658 278822 280894
rect 278266 280338 278502 280574
rect 278586 280338 278822 280574
rect 278266 244658 278502 244894
rect 278586 244658 278822 244894
rect 278266 244338 278502 244574
rect 278586 244338 278822 244574
rect 278266 208658 278502 208894
rect 278586 208658 278822 208894
rect 278266 208338 278502 208574
rect 278586 208338 278822 208574
rect 278266 172658 278502 172894
rect 278586 172658 278822 172894
rect 278266 172338 278502 172574
rect 278586 172338 278822 172574
rect 278266 136658 278502 136894
rect 278586 136658 278822 136894
rect 278266 136338 278502 136574
rect 278586 136338 278822 136574
rect 278266 100658 278502 100894
rect 278586 100658 278822 100894
rect 278266 100338 278502 100574
rect 278586 100338 278822 100574
rect 278266 64658 278502 64894
rect 278586 64658 278822 64894
rect 278266 64338 278502 64574
rect 278586 64338 278822 64574
rect 278266 28658 278502 28894
rect 278586 28658 278822 28894
rect 278266 28338 278502 28574
rect 278586 28338 278822 28574
rect 280826 704602 281062 704838
rect 281146 704602 281382 704838
rect 280826 704282 281062 704518
rect 281146 704282 281382 704518
rect 280826 687218 281062 687454
rect 281146 687218 281382 687454
rect 280826 686898 281062 687134
rect 281146 686898 281382 687134
rect 280826 651218 281062 651454
rect 281146 651218 281382 651454
rect 280826 650898 281062 651134
rect 281146 650898 281382 651134
rect 280826 615218 281062 615454
rect 281146 615218 281382 615454
rect 280826 614898 281062 615134
rect 281146 614898 281382 615134
rect 280826 579218 281062 579454
rect 281146 579218 281382 579454
rect 280826 578898 281062 579134
rect 281146 578898 281382 579134
rect 280826 543218 281062 543454
rect 281146 543218 281382 543454
rect 280826 542898 281062 543134
rect 281146 542898 281382 543134
rect 280826 507218 281062 507454
rect 281146 507218 281382 507454
rect 280826 506898 281062 507134
rect 281146 506898 281382 507134
rect 280826 471218 281062 471454
rect 281146 471218 281382 471454
rect 280826 470898 281062 471134
rect 281146 470898 281382 471134
rect 280826 435218 281062 435454
rect 281146 435218 281382 435454
rect 280826 434898 281062 435134
rect 281146 434898 281382 435134
rect 280826 399218 281062 399454
rect 281146 399218 281382 399454
rect 280826 398898 281062 399134
rect 281146 398898 281382 399134
rect 280826 363218 281062 363454
rect 281146 363218 281382 363454
rect 280826 362898 281062 363134
rect 281146 362898 281382 363134
rect 280826 327218 281062 327454
rect 281146 327218 281382 327454
rect 280826 326898 281062 327134
rect 281146 326898 281382 327134
rect 280826 291218 281062 291454
rect 281146 291218 281382 291454
rect 280826 290898 281062 291134
rect 281146 290898 281382 291134
rect 280826 255218 281062 255454
rect 281146 255218 281382 255454
rect 280826 254898 281062 255134
rect 281146 254898 281382 255134
rect 280826 219218 281062 219454
rect 281146 219218 281382 219454
rect 280826 218898 281062 219134
rect 281146 218898 281382 219134
rect 280826 183218 281062 183454
rect 281146 183218 281382 183454
rect 280826 182898 281062 183134
rect 281146 182898 281382 183134
rect 280826 147218 281062 147454
rect 281146 147218 281382 147454
rect 280826 146898 281062 147134
rect 281146 146898 281382 147134
rect 280826 111218 281062 111454
rect 281146 111218 281382 111454
rect 280826 110898 281062 111134
rect 281146 110898 281382 111134
rect 280826 75218 281062 75454
rect 281146 75218 281382 75454
rect 280826 74898 281062 75134
rect 281146 74898 281382 75134
rect 280826 39218 281062 39454
rect 281146 39218 281382 39454
rect 280826 38898 281062 39134
rect 281146 38898 281382 39134
rect 280826 3218 281062 3454
rect 281146 3218 281382 3454
rect 280826 2898 281062 3134
rect 281146 2898 281382 3134
rect 280826 -582 281062 -346
rect 281146 -582 281382 -346
rect 280826 -902 281062 -666
rect 281146 -902 281382 -666
rect 291986 710362 292222 710598
rect 292306 710362 292542 710598
rect 291986 710042 292222 710278
rect 292306 710042 292542 710278
rect 288266 708442 288502 708678
rect 288586 708442 288822 708678
rect 288266 708122 288502 708358
rect 288586 708122 288822 708358
rect 281986 680378 282222 680614
rect 282306 680378 282542 680614
rect 281986 680058 282222 680294
rect 282306 680058 282542 680294
rect 281986 644378 282222 644614
rect 282306 644378 282542 644614
rect 281986 644058 282222 644294
rect 282306 644058 282542 644294
rect 281986 608378 282222 608614
rect 282306 608378 282542 608614
rect 281986 608058 282222 608294
rect 282306 608058 282542 608294
rect 281986 572378 282222 572614
rect 282306 572378 282542 572614
rect 281986 572058 282222 572294
rect 282306 572058 282542 572294
rect 281986 536378 282222 536614
rect 282306 536378 282542 536614
rect 281986 536058 282222 536294
rect 282306 536058 282542 536294
rect 281986 500378 282222 500614
rect 282306 500378 282542 500614
rect 281986 500058 282222 500294
rect 282306 500058 282542 500294
rect 281986 464378 282222 464614
rect 282306 464378 282542 464614
rect 281986 464058 282222 464294
rect 282306 464058 282542 464294
rect 281986 428378 282222 428614
rect 282306 428378 282542 428614
rect 281986 428058 282222 428294
rect 282306 428058 282542 428294
rect 281986 392378 282222 392614
rect 282306 392378 282542 392614
rect 281986 392058 282222 392294
rect 282306 392058 282542 392294
rect 281986 356378 282222 356614
rect 282306 356378 282542 356614
rect 281986 356058 282222 356294
rect 282306 356058 282542 356294
rect 281986 320378 282222 320614
rect 282306 320378 282542 320614
rect 281986 320058 282222 320294
rect 282306 320058 282542 320294
rect 281986 284378 282222 284614
rect 282306 284378 282542 284614
rect 281986 284058 282222 284294
rect 282306 284058 282542 284294
rect 281986 248378 282222 248614
rect 282306 248378 282542 248614
rect 281986 248058 282222 248294
rect 282306 248058 282542 248294
rect 281986 212378 282222 212614
rect 282306 212378 282542 212614
rect 281986 212058 282222 212294
rect 282306 212058 282542 212294
rect 281986 176378 282222 176614
rect 282306 176378 282542 176614
rect 281986 176058 282222 176294
rect 282306 176058 282542 176294
rect 281986 140378 282222 140614
rect 282306 140378 282542 140614
rect 281986 140058 282222 140294
rect 282306 140058 282542 140294
rect 281986 104378 282222 104614
rect 282306 104378 282542 104614
rect 281986 104058 282222 104294
rect 282306 104058 282542 104294
rect 281986 68378 282222 68614
rect 282306 68378 282542 68614
rect 281986 68058 282222 68294
rect 282306 68058 282542 68294
rect 281986 32378 282222 32614
rect 282306 32378 282542 32614
rect 281986 32058 282222 32294
rect 282306 32058 282542 32294
rect 278266 -5382 278502 -5146
rect 278586 -5382 278822 -5146
rect 278266 -5702 278502 -5466
rect 278586 -5702 278822 -5466
rect 271986 -6342 272222 -6106
rect 272306 -6342 272542 -6106
rect 271986 -6662 272222 -6426
rect 272306 -6662 272542 -6426
rect 284546 706522 284782 706758
rect 284866 706522 285102 706758
rect 284546 706202 284782 706438
rect 284866 706202 285102 706438
rect 284546 690938 284782 691174
rect 284866 690938 285102 691174
rect 284546 690618 284782 690854
rect 284866 690618 285102 690854
rect 284546 654938 284782 655174
rect 284866 654938 285102 655174
rect 284546 654618 284782 654854
rect 284866 654618 285102 654854
rect 284546 618938 284782 619174
rect 284866 618938 285102 619174
rect 284546 618618 284782 618854
rect 284866 618618 285102 618854
rect 284546 582938 284782 583174
rect 284866 582938 285102 583174
rect 284546 582618 284782 582854
rect 284866 582618 285102 582854
rect 284546 546938 284782 547174
rect 284866 546938 285102 547174
rect 284546 546618 284782 546854
rect 284866 546618 285102 546854
rect 284546 510938 284782 511174
rect 284866 510938 285102 511174
rect 284546 510618 284782 510854
rect 284866 510618 285102 510854
rect 284546 474938 284782 475174
rect 284866 474938 285102 475174
rect 284546 474618 284782 474854
rect 284866 474618 285102 474854
rect 284546 438938 284782 439174
rect 284866 438938 285102 439174
rect 284546 438618 284782 438854
rect 284866 438618 285102 438854
rect 284546 402938 284782 403174
rect 284866 402938 285102 403174
rect 284546 402618 284782 402854
rect 284866 402618 285102 402854
rect 284546 366938 284782 367174
rect 284866 366938 285102 367174
rect 284546 366618 284782 366854
rect 284866 366618 285102 366854
rect 284546 330938 284782 331174
rect 284866 330938 285102 331174
rect 284546 330618 284782 330854
rect 284866 330618 285102 330854
rect 284546 294938 284782 295174
rect 284866 294938 285102 295174
rect 284546 294618 284782 294854
rect 284866 294618 285102 294854
rect 284546 258938 284782 259174
rect 284866 258938 285102 259174
rect 284546 258618 284782 258854
rect 284866 258618 285102 258854
rect 284546 222938 284782 223174
rect 284866 222938 285102 223174
rect 284546 222618 284782 222854
rect 284866 222618 285102 222854
rect 284546 186938 284782 187174
rect 284866 186938 285102 187174
rect 284546 186618 284782 186854
rect 284866 186618 285102 186854
rect 284546 150938 284782 151174
rect 284866 150938 285102 151174
rect 284546 150618 284782 150854
rect 284866 150618 285102 150854
rect 284546 114938 284782 115174
rect 284866 114938 285102 115174
rect 284546 114618 284782 114854
rect 284866 114618 285102 114854
rect 284546 78938 284782 79174
rect 284866 78938 285102 79174
rect 284546 78618 284782 78854
rect 284866 78618 285102 78854
rect 284546 42938 284782 43174
rect 284866 42938 285102 43174
rect 284546 42618 284782 42854
rect 284866 42618 285102 42854
rect 284546 6938 284782 7174
rect 284866 6938 285102 7174
rect 284546 6618 284782 6854
rect 284866 6618 285102 6854
rect 284546 -2502 284782 -2266
rect 284866 -2502 285102 -2266
rect 284546 -2822 284782 -2586
rect 284866 -2822 285102 -2586
rect 288266 694658 288502 694894
rect 288586 694658 288822 694894
rect 288266 694338 288502 694574
rect 288586 694338 288822 694574
rect 288266 658658 288502 658894
rect 288586 658658 288822 658894
rect 288266 658338 288502 658574
rect 288586 658338 288822 658574
rect 288266 622658 288502 622894
rect 288586 622658 288822 622894
rect 288266 622338 288502 622574
rect 288586 622338 288822 622574
rect 288266 586658 288502 586894
rect 288586 586658 288822 586894
rect 288266 586338 288502 586574
rect 288586 586338 288822 586574
rect 288266 550658 288502 550894
rect 288586 550658 288822 550894
rect 288266 550338 288502 550574
rect 288586 550338 288822 550574
rect 288266 514658 288502 514894
rect 288586 514658 288822 514894
rect 288266 514338 288502 514574
rect 288586 514338 288822 514574
rect 288266 478658 288502 478894
rect 288586 478658 288822 478894
rect 288266 478338 288502 478574
rect 288586 478338 288822 478574
rect 288266 442658 288502 442894
rect 288586 442658 288822 442894
rect 288266 442338 288502 442574
rect 288586 442338 288822 442574
rect 288266 406658 288502 406894
rect 288586 406658 288822 406894
rect 288266 406338 288502 406574
rect 288586 406338 288822 406574
rect 288266 370658 288502 370894
rect 288586 370658 288822 370894
rect 288266 370338 288502 370574
rect 288586 370338 288822 370574
rect 288266 334658 288502 334894
rect 288586 334658 288822 334894
rect 288266 334338 288502 334574
rect 288586 334338 288822 334574
rect 288266 298658 288502 298894
rect 288586 298658 288822 298894
rect 288266 298338 288502 298574
rect 288586 298338 288822 298574
rect 288266 262658 288502 262894
rect 288586 262658 288822 262894
rect 288266 262338 288502 262574
rect 288586 262338 288822 262574
rect 288266 226658 288502 226894
rect 288586 226658 288822 226894
rect 288266 226338 288502 226574
rect 288586 226338 288822 226574
rect 288266 190658 288502 190894
rect 288586 190658 288822 190894
rect 288266 190338 288502 190574
rect 288586 190338 288822 190574
rect 288266 154658 288502 154894
rect 288586 154658 288822 154894
rect 288266 154338 288502 154574
rect 288586 154338 288822 154574
rect 288266 118658 288502 118894
rect 288586 118658 288822 118894
rect 288266 118338 288502 118574
rect 288586 118338 288822 118574
rect 288266 82658 288502 82894
rect 288586 82658 288822 82894
rect 288266 82338 288502 82574
rect 288586 82338 288822 82574
rect 288266 46658 288502 46894
rect 288586 46658 288822 46894
rect 288266 46338 288502 46574
rect 288586 46338 288822 46574
rect 288266 10658 288502 10894
rect 288586 10658 288822 10894
rect 288266 10338 288502 10574
rect 288586 10338 288822 10574
rect 290826 705562 291062 705798
rect 291146 705562 291382 705798
rect 290826 705242 291062 705478
rect 291146 705242 291382 705478
rect 290826 669218 291062 669454
rect 291146 669218 291382 669454
rect 290826 668898 291062 669134
rect 291146 668898 291382 669134
rect 290826 633218 291062 633454
rect 291146 633218 291382 633454
rect 290826 632898 291062 633134
rect 291146 632898 291382 633134
rect 290826 597218 291062 597454
rect 291146 597218 291382 597454
rect 290826 596898 291062 597134
rect 291146 596898 291382 597134
rect 290826 561218 291062 561454
rect 291146 561218 291382 561454
rect 290826 560898 291062 561134
rect 291146 560898 291382 561134
rect 290826 525218 291062 525454
rect 291146 525218 291382 525454
rect 290826 524898 291062 525134
rect 291146 524898 291382 525134
rect 290826 489218 291062 489454
rect 291146 489218 291382 489454
rect 290826 488898 291062 489134
rect 291146 488898 291382 489134
rect 290826 453218 291062 453454
rect 291146 453218 291382 453454
rect 290826 452898 291062 453134
rect 291146 452898 291382 453134
rect 290826 417218 291062 417454
rect 291146 417218 291382 417454
rect 290826 416898 291062 417134
rect 291146 416898 291382 417134
rect 290826 381218 291062 381454
rect 291146 381218 291382 381454
rect 290826 380898 291062 381134
rect 291146 380898 291382 381134
rect 290826 345218 291062 345454
rect 291146 345218 291382 345454
rect 290826 344898 291062 345134
rect 291146 344898 291382 345134
rect 290826 309218 291062 309454
rect 291146 309218 291382 309454
rect 290826 308898 291062 309134
rect 291146 308898 291382 309134
rect 290826 273218 291062 273454
rect 291146 273218 291382 273454
rect 290826 272898 291062 273134
rect 291146 272898 291382 273134
rect 290826 237218 291062 237454
rect 291146 237218 291382 237454
rect 290826 236898 291062 237134
rect 291146 236898 291382 237134
rect 290826 201218 291062 201454
rect 291146 201218 291382 201454
rect 290826 200898 291062 201134
rect 291146 200898 291382 201134
rect 290826 165218 291062 165454
rect 291146 165218 291382 165454
rect 290826 164898 291062 165134
rect 291146 164898 291382 165134
rect 290826 129218 291062 129454
rect 291146 129218 291382 129454
rect 290826 128898 291062 129134
rect 291146 128898 291382 129134
rect 290826 93218 291062 93454
rect 291146 93218 291382 93454
rect 290826 92898 291062 93134
rect 291146 92898 291382 93134
rect 290826 57218 291062 57454
rect 291146 57218 291382 57454
rect 290826 56898 291062 57134
rect 291146 56898 291382 57134
rect 290826 21218 291062 21454
rect 291146 21218 291382 21454
rect 290826 20898 291062 21134
rect 291146 20898 291382 21134
rect 290826 -1542 291062 -1306
rect 291146 -1542 291382 -1306
rect 290826 -1862 291062 -1626
rect 291146 -1862 291382 -1626
rect 301986 711322 302222 711558
rect 302306 711322 302542 711558
rect 301986 711002 302222 711238
rect 302306 711002 302542 711238
rect 298266 709402 298502 709638
rect 298586 709402 298822 709638
rect 298266 709082 298502 709318
rect 298586 709082 298822 709318
rect 291986 698378 292222 698614
rect 292306 698378 292542 698614
rect 291986 698058 292222 698294
rect 292306 698058 292542 698294
rect 291986 662378 292222 662614
rect 292306 662378 292542 662614
rect 291986 662058 292222 662294
rect 292306 662058 292542 662294
rect 291986 626378 292222 626614
rect 292306 626378 292542 626614
rect 291986 626058 292222 626294
rect 292306 626058 292542 626294
rect 291986 590378 292222 590614
rect 292306 590378 292542 590614
rect 291986 590058 292222 590294
rect 292306 590058 292542 590294
rect 291986 554378 292222 554614
rect 292306 554378 292542 554614
rect 291986 554058 292222 554294
rect 292306 554058 292542 554294
rect 291986 518378 292222 518614
rect 292306 518378 292542 518614
rect 291986 518058 292222 518294
rect 292306 518058 292542 518294
rect 291986 482378 292222 482614
rect 292306 482378 292542 482614
rect 291986 482058 292222 482294
rect 292306 482058 292542 482294
rect 291986 446378 292222 446614
rect 292306 446378 292542 446614
rect 291986 446058 292222 446294
rect 292306 446058 292542 446294
rect 291986 410378 292222 410614
rect 292306 410378 292542 410614
rect 291986 410058 292222 410294
rect 292306 410058 292542 410294
rect 291986 374378 292222 374614
rect 292306 374378 292542 374614
rect 291986 374058 292222 374294
rect 292306 374058 292542 374294
rect 291986 338378 292222 338614
rect 292306 338378 292542 338614
rect 291986 338058 292222 338294
rect 292306 338058 292542 338294
rect 291986 302378 292222 302614
rect 292306 302378 292542 302614
rect 291986 302058 292222 302294
rect 292306 302058 292542 302294
rect 291986 266378 292222 266614
rect 292306 266378 292542 266614
rect 291986 266058 292222 266294
rect 292306 266058 292542 266294
rect 291986 230378 292222 230614
rect 292306 230378 292542 230614
rect 291986 230058 292222 230294
rect 292306 230058 292542 230294
rect 291986 194378 292222 194614
rect 292306 194378 292542 194614
rect 291986 194058 292222 194294
rect 292306 194058 292542 194294
rect 291986 158378 292222 158614
rect 292306 158378 292542 158614
rect 291986 158058 292222 158294
rect 292306 158058 292542 158294
rect 291986 122378 292222 122614
rect 292306 122378 292542 122614
rect 291986 122058 292222 122294
rect 292306 122058 292542 122294
rect 291986 86378 292222 86614
rect 292306 86378 292542 86614
rect 291986 86058 292222 86294
rect 292306 86058 292542 86294
rect 291986 50378 292222 50614
rect 292306 50378 292542 50614
rect 291986 50058 292222 50294
rect 292306 50058 292542 50294
rect 291986 14378 292222 14614
rect 292306 14378 292542 14614
rect 291986 14058 292222 14294
rect 292306 14058 292542 14294
rect 288266 -4422 288502 -4186
rect 288586 -4422 288822 -4186
rect 288266 -4742 288502 -4506
rect 288586 -4742 288822 -4506
rect 281986 -7302 282222 -7066
rect 282306 -7302 282542 -7066
rect 281986 -7622 282222 -7386
rect 282306 -7622 282542 -7386
rect 294546 707482 294782 707718
rect 294866 707482 295102 707718
rect 294546 707162 294782 707398
rect 294866 707162 295102 707398
rect 294546 672938 294782 673174
rect 294866 672938 295102 673174
rect 294546 672618 294782 672854
rect 294866 672618 295102 672854
rect 294546 636938 294782 637174
rect 294866 636938 295102 637174
rect 294546 636618 294782 636854
rect 294866 636618 295102 636854
rect 294546 600938 294782 601174
rect 294866 600938 295102 601174
rect 294546 600618 294782 600854
rect 294866 600618 295102 600854
rect 294546 564938 294782 565174
rect 294866 564938 295102 565174
rect 294546 564618 294782 564854
rect 294866 564618 295102 564854
rect 294546 528938 294782 529174
rect 294866 528938 295102 529174
rect 294546 528618 294782 528854
rect 294866 528618 295102 528854
rect 294546 492938 294782 493174
rect 294866 492938 295102 493174
rect 294546 492618 294782 492854
rect 294866 492618 295102 492854
rect 294546 456938 294782 457174
rect 294866 456938 295102 457174
rect 294546 456618 294782 456854
rect 294866 456618 295102 456854
rect 294546 420938 294782 421174
rect 294866 420938 295102 421174
rect 294546 420618 294782 420854
rect 294866 420618 295102 420854
rect 294546 384938 294782 385174
rect 294866 384938 295102 385174
rect 294546 384618 294782 384854
rect 294866 384618 295102 384854
rect 294546 348938 294782 349174
rect 294866 348938 295102 349174
rect 294546 348618 294782 348854
rect 294866 348618 295102 348854
rect 294546 312938 294782 313174
rect 294866 312938 295102 313174
rect 294546 312618 294782 312854
rect 294866 312618 295102 312854
rect 294546 276938 294782 277174
rect 294866 276938 295102 277174
rect 294546 276618 294782 276854
rect 294866 276618 295102 276854
rect 294546 240938 294782 241174
rect 294866 240938 295102 241174
rect 294546 240618 294782 240854
rect 294866 240618 295102 240854
rect 294546 204938 294782 205174
rect 294866 204938 295102 205174
rect 294546 204618 294782 204854
rect 294866 204618 295102 204854
rect 294546 168938 294782 169174
rect 294866 168938 295102 169174
rect 294546 168618 294782 168854
rect 294866 168618 295102 168854
rect 294546 132938 294782 133174
rect 294866 132938 295102 133174
rect 294546 132618 294782 132854
rect 294866 132618 295102 132854
rect 294546 96938 294782 97174
rect 294866 96938 295102 97174
rect 294546 96618 294782 96854
rect 294866 96618 295102 96854
rect 294546 60938 294782 61174
rect 294866 60938 295102 61174
rect 294546 60618 294782 60854
rect 294866 60618 295102 60854
rect 294546 24938 294782 25174
rect 294866 24938 295102 25174
rect 294546 24618 294782 24854
rect 294866 24618 295102 24854
rect 294546 -3462 294782 -3226
rect 294866 -3462 295102 -3226
rect 294546 -3782 294782 -3546
rect 294866 -3782 295102 -3546
rect 298266 676658 298502 676894
rect 298586 676658 298822 676894
rect 298266 676338 298502 676574
rect 298586 676338 298822 676574
rect 298266 640658 298502 640894
rect 298586 640658 298822 640894
rect 298266 640338 298502 640574
rect 298586 640338 298822 640574
rect 298266 604658 298502 604894
rect 298586 604658 298822 604894
rect 298266 604338 298502 604574
rect 298586 604338 298822 604574
rect 298266 568658 298502 568894
rect 298586 568658 298822 568894
rect 298266 568338 298502 568574
rect 298586 568338 298822 568574
rect 298266 532658 298502 532894
rect 298586 532658 298822 532894
rect 298266 532338 298502 532574
rect 298586 532338 298822 532574
rect 298266 496658 298502 496894
rect 298586 496658 298822 496894
rect 298266 496338 298502 496574
rect 298586 496338 298822 496574
rect 298266 460658 298502 460894
rect 298586 460658 298822 460894
rect 298266 460338 298502 460574
rect 298586 460338 298822 460574
rect 298266 424658 298502 424894
rect 298586 424658 298822 424894
rect 298266 424338 298502 424574
rect 298586 424338 298822 424574
rect 298266 388658 298502 388894
rect 298586 388658 298822 388894
rect 298266 388338 298502 388574
rect 298586 388338 298822 388574
rect 298266 352658 298502 352894
rect 298586 352658 298822 352894
rect 298266 352338 298502 352574
rect 298586 352338 298822 352574
rect 298266 316658 298502 316894
rect 298586 316658 298822 316894
rect 298266 316338 298502 316574
rect 298586 316338 298822 316574
rect 298266 280658 298502 280894
rect 298586 280658 298822 280894
rect 298266 280338 298502 280574
rect 298586 280338 298822 280574
rect 298266 244658 298502 244894
rect 298586 244658 298822 244894
rect 298266 244338 298502 244574
rect 298586 244338 298822 244574
rect 298266 208658 298502 208894
rect 298586 208658 298822 208894
rect 298266 208338 298502 208574
rect 298586 208338 298822 208574
rect 298266 172658 298502 172894
rect 298586 172658 298822 172894
rect 298266 172338 298502 172574
rect 298586 172338 298822 172574
rect 298266 136658 298502 136894
rect 298586 136658 298822 136894
rect 298266 136338 298502 136574
rect 298586 136338 298822 136574
rect 298266 100658 298502 100894
rect 298586 100658 298822 100894
rect 298266 100338 298502 100574
rect 298586 100338 298822 100574
rect 298266 64658 298502 64894
rect 298586 64658 298822 64894
rect 298266 64338 298502 64574
rect 298586 64338 298822 64574
rect 298266 28658 298502 28894
rect 298586 28658 298822 28894
rect 298266 28338 298502 28574
rect 298586 28338 298822 28574
rect 300826 704602 301062 704838
rect 301146 704602 301382 704838
rect 300826 704282 301062 704518
rect 301146 704282 301382 704518
rect 300826 687218 301062 687454
rect 301146 687218 301382 687454
rect 300826 686898 301062 687134
rect 301146 686898 301382 687134
rect 300826 651218 301062 651454
rect 301146 651218 301382 651454
rect 300826 650898 301062 651134
rect 301146 650898 301382 651134
rect 300826 615218 301062 615454
rect 301146 615218 301382 615454
rect 300826 614898 301062 615134
rect 301146 614898 301382 615134
rect 300826 579218 301062 579454
rect 301146 579218 301382 579454
rect 300826 578898 301062 579134
rect 301146 578898 301382 579134
rect 300826 543218 301062 543454
rect 301146 543218 301382 543454
rect 300826 542898 301062 543134
rect 301146 542898 301382 543134
rect 300826 507218 301062 507454
rect 301146 507218 301382 507454
rect 300826 506898 301062 507134
rect 301146 506898 301382 507134
rect 300826 471218 301062 471454
rect 301146 471218 301382 471454
rect 300826 470898 301062 471134
rect 301146 470898 301382 471134
rect 300826 435218 301062 435454
rect 301146 435218 301382 435454
rect 300826 434898 301062 435134
rect 301146 434898 301382 435134
rect 300826 399218 301062 399454
rect 301146 399218 301382 399454
rect 300826 398898 301062 399134
rect 301146 398898 301382 399134
rect 300826 363218 301062 363454
rect 301146 363218 301382 363454
rect 300826 362898 301062 363134
rect 301146 362898 301382 363134
rect 300826 327218 301062 327454
rect 301146 327218 301382 327454
rect 300826 326898 301062 327134
rect 301146 326898 301382 327134
rect 300826 291218 301062 291454
rect 301146 291218 301382 291454
rect 300826 290898 301062 291134
rect 301146 290898 301382 291134
rect 300826 255218 301062 255454
rect 301146 255218 301382 255454
rect 300826 254898 301062 255134
rect 301146 254898 301382 255134
rect 300826 219218 301062 219454
rect 301146 219218 301382 219454
rect 300826 218898 301062 219134
rect 301146 218898 301382 219134
rect 300826 183218 301062 183454
rect 301146 183218 301382 183454
rect 300826 182898 301062 183134
rect 301146 182898 301382 183134
rect 300826 147218 301062 147454
rect 301146 147218 301382 147454
rect 300826 146898 301062 147134
rect 301146 146898 301382 147134
rect 300826 111218 301062 111454
rect 301146 111218 301382 111454
rect 300826 110898 301062 111134
rect 301146 110898 301382 111134
rect 300826 75218 301062 75454
rect 301146 75218 301382 75454
rect 300826 74898 301062 75134
rect 301146 74898 301382 75134
rect 300826 39218 301062 39454
rect 301146 39218 301382 39454
rect 300826 38898 301062 39134
rect 301146 38898 301382 39134
rect 300826 3218 301062 3454
rect 301146 3218 301382 3454
rect 300826 2898 301062 3134
rect 301146 2898 301382 3134
rect 300826 -582 301062 -346
rect 301146 -582 301382 -346
rect 300826 -902 301062 -666
rect 301146 -902 301382 -666
rect 311986 710362 312222 710598
rect 312306 710362 312542 710598
rect 311986 710042 312222 710278
rect 312306 710042 312542 710278
rect 308266 708442 308502 708678
rect 308586 708442 308822 708678
rect 308266 708122 308502 708358
rect 308586 708122 308822 708358
rect 301986 680378 302222 680614
rect 302306 680378 302542 680614
rect 301986 680058 302222 680294
rect 302306 680058 302542 680294
rect 301986 644378 302222 644614
rect 302306 644378 302542 644614
rect 301986 644058 302222 644294
rect 302306 644058 302542 644294
rect 301986 608378 302222 608614
rect 302306 608378 302542 608614
rect 301986 608058 302222 608294
rect 302306 608058 302542 608294
rect 301986 572378 302222 572614
rect 302306 572378 302542 572614
rect 301986 572058 302222 572294
rect 302306 572058 302542 572294
rect 301986 536378 302222 536614
rect 302306 536378 302542 536614
rect 301986 536058 302222 536294
rect 302306 536058 302542 536294
rect 301986 500378 302222 500614
rect 302306 500378 302542 500614
rect 301986 500058 302222 500294
rect 302306 500058 302542 500294
rect 301986 464378 302222 464614
rect 302306 464378 302542 464614
rect 301986 464058 302222 464294
rect 302306 464058 302542 464294
rect 301986 428378 302222 428614
rect 302306 428378 302542 428614
rect 301986 428058 302222 428294
rect 302306 428058 302542 428294
rect 301986 392378 302222 392614
rect 302306 392378 302542 392614
rect 301986 392058 302222 392294
rect 302306 392058 302542 392294
rect 301986 356378 302222 356614
rect 302306 356378 302542 356614
rect 301986 356058 302222 356294
rect 302306 356058 302542 356294
rect 301986 320378 302222 320614
rect 302306 320378 302542 320614
rect 301986 320058 302222 320294
rect 302306 320058 302542 320294
rect 301986 284378 302222 284614
rect 302306 284378 302542 284614
rect 301986 284058 302222 284294
rect 302306 284058 302542 284294
rect 301986 248378 302222 248614
rect 302306 248378 302542 248614
rect 301986 248058 302222 248294
rect 302306 248058 302542 248294
rect 301986 212378 302222 212614
rect 302306 212378 302542 212614
rect 301986 212058 302222 212294
rect 302306 212058 302542 212294
rect 301986 176378 302222 176614
rect 302306 176378 302542 176614
rect 301986 176058 302222 176294
rect 302306 176058 302542 176294
rect 301986 140378 302222 140614
rect 302306 140378 302542 140614
rect 301986 140058 302222 140294
rect 302306 140058 302542 140294
rect 301986 104378 302222 104614
rect 302306 104378 302542 104614
rect 301986 104058 302222 104294
rect 302306 104058 302542 104294
rect 301986 68378 302222 68614
rect 302306 68378 302542 68614
rect 301986 68058 302222 68294
rect 302306 68058 302542 68294
rect 301986 32378 302222 32614
rect 302306 32378 302542 32614
rect 301986 32058 302222 32294
rect 302306 32058 302542 32294
rect 298266 -5382 298502 -5146
rect 298586 -5382 298822 -5146
rect 298266 -5702 298502 -5466
rect 298586 -5702 298822 -5466
rect 291986 -6342 292222 -6106
rect 292306 -6342 292542 -6106
rect 291986 -6662 292222 -6426
rect 292306 -6662 292542 -6426
rect 304546 706522 304782 706758
rect 304866 706522 305102 706758
rect 304546 706202 304782 706438
rect 304866 706202 305102 706438
rect 304546 690938 304782 691174
rect 304866 690938 305102 691174
rect 304546 690618 304782 690854
rect 304866 690618 305102 690854
rect 304546 654938 304782 655174
rect 304866 654938 305102 655174
rect 304546 654618 304782 654854
rect 304866 654618 305102 654854
rect 304546 618938 304782 619174
rect 304866 618938 305102 619174
rect 304546 618618 304782 618854
rect 304866 618618 305102 618854
rect 304546 582938 304782 583174
rect 304866 582938 305102 583174
rect 304546 582618 304782 582854
rect 304866 582618 305102 582854
rect 304546 546938 304782 547174
rect 304866 546938 305102 547174
rect 304546 546618 304782 546854
rect 304866 546618 305102 546854
rect 304546 510938 304782 511174
rect 304866 510938 305102 511174
rect 304546 510618 304782 510854
rect 304866 510618 305102 510854
rect 304546 474938 304782 475174
rect 304866 474938 305102 475174
rect 304546 474618 304782 474854
rect 304866 474618 305102 474854
rect 304546 438938 304782 439174
rect 304866 438938 305102 439174
rect 304546 438618 304782 438854
rect 304866 438618 305102 438854
rect 304546 402938 304782 403174
rect 304866 402938 305102 403174
rect 304546 402618 304782 402854
rect 304866 402618 305102 402854
rect 304546 366938 304782 367174
rect 304866 366938 305102 367174
rect 304546 366618 304782 366854
rect 304866 366618 305102 366854
rect 304546 330938 304782 331174
rect 304866 330938 305102 331174
rect 304546 330618 304782 330854
rect 304866 330618 305102 330854
rect 304546 294938 304782 295174
rect 304866 294938 305102 295174
rect 304546 294618 304782 294854
rect 304866 294618 305102 294854
rect 304546 258938 304782 259174
rect 304866 258938 305102 259174
rect 304546 258618 304782 258854
rect 304866 258618 305102 258854
rect 304546 222938 304782 223174
rect 304866 222938 305102 223174
rect 304546 222618 304782 222854
rect 304866 222618 305102 222854
rect 304546 186938 304782 187174
rect 304866 186938 305102 187174
rect 304546 186618 304782 186854
rect 304866 186618 305102 186854
rect 304546 150938 304782 151174
rect 304866 150938 305102 151174
rect 304546 150618 304782 150854
rect 304866 150618 305102 150854
rect 304546 114938 304782 115174
rect 304866 114938 305102 115174
rect 304546 114618 304782 114854
rect 304866 114618 305102 114854
rect 304546 78938 304782 79174
rect 304866 78938 305102 79174
rect 304546 78618 304782 78854
rect 304866 78618 305102 78854
rect 304546 42938 304782 43174
rect 304866 42938 305102 43174
rect 304546 42618 304782 42854
rect 304866 42618 305102 42854
rect 304546 6938 304782 7174
rect 304866 6938 305102 7174
rect 304546 6618 304782 6854
rect 304866 6618 305102 6854
rect 304546 -2502 304782 -2266
rect 304866 -2502 305102 -2266
rect 304546 -2822 304782 -2586
rect 304866 -2822 305102 -2586
rect 308266 694658 308502 694894
rect 308586 694658 308822 694894
rect 308266 694338 308502 694574
rect 308586 694338 308822 694574
rect 308266 658658 308502 658894
rect 308586 658658 308822 658894
rect 308266 658338 308502 658574
rect 308586 658338 308822 658574
rect 308266 622658 308502 622894
rect 308586 622658 308822 622894
rect 308266 622338 308502 622574
rect 308586 622338 308822 622574
rect 308266 586658 308502 586894
rect 308586 586658 308822 586894
rect 308266 586338 308502 586574
rect 308586 586338 308822 586574
rect 308266 550658 308502 550894
rect 308586 550658 308822 550894
rect 308266 550338 308502 550574
rect 308586 550338 308822 550574
rect 308266 514658 308502 514894
rect 308586 514658 308822 514894
rect 308266 514338 308502 514574
rect 308586 514338 308822 514574
rect 308266 478658 308502 478894
rect 308586 478658 308822 478894
rect 308266 478338 308502 478574
rect 308586 478338 308822 478574
rect 308266 442658 308502 442894
rect 308586 442658 308822 442894
rect 308266 442338 308502 442574
rect 308586 442338 308822 442574
rect 308266 406658 308502 406894
rect 308586 406658 308822 406894
rect 308266 406338 308502 406574
rect 308586 406338 308822 406574
rect 308266 370658 308502 370894
rect 308586 370658 308822 370894
rect 308266 370338 308502 370574
rect 308586 370338 308822 370574
rect 308266 334658 308502 334894
rect 308586 334658 308822 334894
rect 308266 334338 308502 334574
rect 308586 334338 308822 334574
rect 308266 298658 308502 298894
rect 308586 298658 308822 298894
rect 308266 298338 308502 298574
rect 308586 298338 308822 298574
rect 308266 262658 308502 262894
rect 308586 262658 308822 262894
rect 308266 262338 308502 262574
rect 308586 262338 308822 262574
rect 308266 226658 308502 226894
rect 308586 226658 308822 226894
rect 308266 226338 308502 226574
rect 308586 226338 308822 226574
rect 308266 190658 308502 190894
rect 308586 190658 308822 190894
rect 308266 190338 308502 190574
rect 308586 190338 308822 190574
rect 308266 154658 308502 154894
rect 308586 154658 308822 154894
rect 308266 154338 308502 154574
rect 308586 154338 308822 154574
rect 308266 118658 308502 118894
rect 308586 118658 308822 118894
rect 308266 118338 308502 118574
rect 308586 118338 308822 118574
rect 308266 82658 308502 82894
rect 308586 82658 308822 82894
rect 308266 82338 308502 82574
rect 308586 82338 308822 82574
rect 308266 46658 308502 46894
rect 308586 46658 308822 46894
rect 308266 46338 308502 46574
rect 308586 46338 308822 46574
rect 308266 10658 308502 10894
rect 308586 10658 308822 10894
rect 308266 10338 308502 10574
rect 308586 10338 308822 10574
rect 310826 705562 311062 705798
rect 311146 705562 311382 705798
rect 310826 705242 311062 705478
rect 311146 705242 311382 705478
rect 310826 669218 311062 669454
rect 311146 669218 311382 669454
rect 310826 668898 311062 669134
rect 311146 668898 311382 669134
rect 310826 633218 311062 633454
rect 311146 633218 311382 633454
rect 310826 632898 311062 633134
rect 311146 632898 311382 633134
rect 310826 597218 311062 597454
rect 311146 597218 311382 597454
rect 310826 596898 311062 597134
rect 311146 596898 311382 597134
rect 310826 561218 311062 561454
rect 311146 561218 311382 561454
rect 310826 560898 311062 561134
rect 311146 560898 311382 561134
rect 310826 525218 311062 525454
rect 311146 525218 311382 525454
rect 310826 524898 311062 525134
rect 311146 524898 311382 525134
rect 310826 489218 311062 489454
rect 311146 489218 311382 489454
rect 310826 488898 311062 489134
rect 311146 488898 311382 489134
rect 310826 453218 311062 453454
rect 311146 453218 311382 453454
rect 310826 452898 311062 453134
rect 311146 452898 311382 453134
rect 310826 417218 311062 417454
rect 311146 417218 311382 417454
rect 310826 416898 311062 417134
rect 311146 416898 311382 417134
rect 310826 381218 311062 381454
rect 311146 381218 311382 381454
rect 310826 380898 311062 381134
rect 311146 380898 311382 381134
rect 310826 345218 311062 345454
rect 311146 345218 311382 345454
rect 310826 344898 311062 345134
rect 311146 344898 311382 345134
rect 310826 309218 311062 309454
rect 311146 309218 311382 309454
rect 310826 308898 311062 309134
rect 311146 308898 311382 309134
rect 310826 273218 311062 273454
rect 311146 273218 311382 273454
rect 310826 272898 311062 273134
rect 311146 272898 311382 273134
rect 310826 237218 311062 237454
rect 311146 237218 311382 237454
rect 310826 236898 311062 237134
rect 311146 236898 311382 237134
rect 310826 201218 311062 201454
rect 311146 201218 311382 201454
rect 310826 200898 311062 201134
rect 311146 200898 311382 201134
rect 310826 165218 311062 165454
rect 311146 165218 311382 165454
rect 310826 164898 311062 165134
rect 311146 164898 311382 165134
rect 310826 129218 311062 129454
rect 311146 129218 311382 129454
rect 310826 128898 311062 129134
rect 311146 128898 311382 129134
rect 310826 93218 311062 93454
rect 311146 93218 311382 93454
rect 310826 92898 311062 93134
rect 311146 92898 311382 93134
rect 310826 57218 311062 57454
rect 311146 57218 311382 57454
rect 310826 56898 311062 57134
rect 311146 56898 311382 57134
rect 310826 21218 311062 21454
rect 311146 21218 311382 21454
rect 310826 20898 311062 21134
rect 311146 20898 311382 21134
rect 310826 -1542 311062 -1306
rect 311146 -1542 311382 -1306
rect 310826 -1862 311062 -1626
rect 311146 -1862 311382 -1626
rect 321986 711322 322222 711558
rect 322306 711322 322542 711558
rect 321986 711002 322222 711238
rect 322306 711002 322542 711238
rect 318266 709402 318502 709638
rect 318586 709402 318822 709638
rect 318266 709082 318502 709318
rect 318586 709082 318822 709318
rect 311986 698378 312222 698614
rect 312306 698378 312542 698614
rect 311986 698058 312222 698294
rect 312306 698058 312542 698294
rect 311986 662378 312222 662614
rect 312306 662378 312542 662614
rect 311986 662058 312222 662294
rect 312306 662058 312542 662294
rect 311986 626378 312222 626614
rect 312306 626378 312542 626614
rect 311986 626058 312222 626294
rect 312306 626058 312542 626294
rect 311986 590378 312222 590614
rect 312306 590378 312542 590614
rect 311986 590058 312222 590294
rect 312306 590058 312542 590294
rect 311986 554378 312222 554614
rect 312306 554378 312542 554614
rect 311986 554058 312222 554294
rect 312306 554058 312542 554294
rect 311986 518378 312222 518614
rect 312306 518378 312542 518614
rect 311986 518058 312222 518294
rect 312306 518058 312542 518294
rect 311986 482378 312222 482614
rect 312306 482378 312542 482614
rect 311986 482058 312222 482294
rect 312306 482058 312542 482294
rect 311986 446378 312222 446614
rect 312306 446378 312542 446614
rect 311986 446058 312222 446294
rect 312306 446058 312542 446294
rect 311986 410378 312222 410614
rect 312306 410378 312542 410614
rect 311986 410058 312222 410294
rect 312306 410058 312542 410294
rect 311986 374378 312222 374614
rect 312306 374378 312542 374614
rect 311986 374058 312222 374294
rect 312306 374058 312542 374294
rect 311986 338378 312222 338614
rect 312306 338378 312542 338614
rect 311986 338058 312222 338294
rect 312306 338058 312542 338294
rect 311986 302378 312222 302614
rect 312306 302378 312542 302614
rect 311986 302058 312222 302294
rect 312306 302058 312542 302294
rect 311986 266378 312222 266614
rect 312306 266378 312542 266614
rect 311986 266058 312222 266294
rect 312306 266058 312542 266294
rect 311986 230378 312222 230614
rect 312306 230378 312542 230614
rect 311986 230058 312222 230294
rect 312306 230058 312542 230294
rect 311986 194378 312222 194614
rect 312306 194378 312542 194614
rect 311986 194058 312222 194294
rect 312306 194058 312542 194294
rect 311986 158378 312222 158614
rect 312306 158378 312542 158614
rect 311986 158058 312222 158294
rect 312306 158058 312542 158294
rect 311986 122378 312222 122614
rect 312306 122378 312542 122614
rect 311986 122058 312222 122294
rect 312306 122058 312542 122294
rect 311986 86378 312222 86614
rect 312306 86378 312542 86614
rect 311986 86058 312222 86294
rect 312306 86058 312542 86294
rect 311986 50378 312222 50614
rect 312306 50378 312542 50614
rect 311986 50058 312222 50294
rect 312306 50058 312542 50294
rect 311986 14378 312222 14614
rect 312306 14378 312542 14614
rect 311986 14058 312222 14294
rect 312306 14058 312542 14294
rect 308266 -4422 308502 -4186
rect 308586 -4422 308822 -4186
rect 308266 -4742 308502 -4506
rect 308586 -4742 308822 -4506
rect 301986 -7302 302222 -7066
rect 302306 -7302 302542 -7066
rect 301986 -7622 302222 -7386
rect 302306 -7622 302542 -7386
rect 314546 707482 314782 707718
rect 314866 707482 315102 707718
rect 314546 707162 314782 707398
rect 314866 707162 315102 707398
rect 314546 672938 314782 673174
rect 314866 672938 315102 673174
rect 314546 672618 314782 672854
rect 314866 672618 315102 672854
rect 314546 636938 314782 637174
rect 314866 636938 315102 637174
rect 314546 636618 314782 636854
rect 314866 636618 315102 636854
rect 314546 600938 314782 601174
rect 314866 600938 315102 601174
rect 314546 600618 314782 600854
rect 314866 600618 315102 600854
rect 314546 564938 314782 565174
rect 314866 564938 315102 565174
rect 314546 564618 314782 564854
rect 314866 564618 315102 564854
rect 314546 528938 314782 529174
rect 314866 528938 315102 529174
rect 314546 528618 314782 528854
rect 314866 528618 315102 528854
rect 314546 492938 314782 493174
rect 314866 492938 315102 493174
rect 314546 492618 314782 492854
rect 314866 492618 315102 492854
rect 314546 456938 314782 457174
rect 314866 456938 315102 457174
rect 314546 456618 314782 456854
rect 314866 456618 315102 456854
rect 314546 420938 314782 421174
rect 314866 420938 315102 421174
rect 314546 420618 314782 420854
rect 314866 420618 315102 420854
rect 314546 384938 314782 385174
rect 314866 384938 315102 385174
rect 314546 384618 314782 384854
rect 314866 384618 315102 384854
rect 314546 348938 314782 349174
rect 314866 348938 315102 349174
rect 314546 348618 314782 348854
rect 314866 348618 315102 348854
rect 314546 312938 314782 313174
rect 314866 312938 315102 313174
rect 314546 312618 314782 312854
rect 314866 312618 315102 312854
rect 314546 276938 314782 277174
rect 314866 276938 315102 277174
rect 314546 276618 314782 276854
rect 314866 276618 315102 276854
rect 314546 240938 314782 241174
rect 314866 240938 315102 241174
rect 314546 240618 314782 240854
rect 314866 240618 315102 240854
rect 314546 204938 314782 205174
rect 314866 204938 315102 205174
rect 314546 204618 314782 204854
rect 314866 204618 315102 204854
rect 314546 168938 314782 169174
rect 314866 168938 315102 169174
rect 314546 168618 314782 168854
rect 314866 168618 315102 168854
rect 314546 132938 314782 133174
rect 314866 132938 315102 133174
rect 314546 132618 314782 132854
rect 314866 132618 315102 132854
rect 314546 96938 314782 97174
rect 314866 96938 315102 97174
rect 314546 96618 314782 96854
rect 314866 96618 315102 96854
rect 314546 60938 314782 61174
rect 314866 60938 315102 61174
rect 314546 60618 314782 60854
rect 314866 60618 315102 60854
rect 314546 24938 314782 25174
rect 314866 24938 315102 25174
rect 314546 24618 314782 24854
rect 314866 24618 315102 24854
rect 314546 -3462 314782 -3226
rect 314866 -3462 315102 -3226
rect 314546 -3782 314782 -3546
rect 314866 -3782 315102 -3546
rect 318266 676658 318502 676894
rect 318586 676658 318822 676894
rect 318266 676338 318502 676574
rect 318586 676338 318822 676574
rect 318266 640658 318502 640894
rect 318586 640658 318822 640894
rect 318266 640338 318502 640574
rect 318586 640338 318822 640574
rect 318266 604658 318502 604894
rect 318586 604658 318822 604894
rect 318266 604338 318502 604574
rect 318586 604338 318822 604574
rect 318266 568658 318502 568894
rect 318586 568658 318822 568894
rect 318266 568338 318502 568574
rect 318586 568338 318822 568574
rect 318266 532658 318502 532894
rect 318586 532658 318822 532894
rect 318266 532338 318502 532574
rect 318586 532338 318822 532574
rect 318266 496658 318502 496894
rect 318586 496658 318822 496894
rect 318266 496338 318502 496574
rect 318586 496338 318822 496574
rect 318266 460658 318502 460894
rect 318586 460658 318822 460894
rect 318266 460338 318502 460574
rect 318586 460338 318822 460574
rect 318266 424658 318502 424894
rect 318586 424658 318822 424894
rect 318266 424338 318502 424574
rect 318586 424338 318822 424574
rect 318266 388658 318502 388894
rect 318586 388658 318822 388894
rect 318266 388338 318502 388574
rect 318586 388338 318822 388574
rect 318266 352658 318502 352894
rect 318586 352658 318822 352894
rect 318266 352338 318502 352574
rect 318586 352338 318822 352574
rect 318266 316658 318502 316894
rect 318586 316658 318822 316894
rect 318266 316338 318502 316574
rect 318586 316338 318822 316574
rect 318266 280658 318502 280894
rect 318586 280658 318822 280894
rect 318266 280338 318502 280574
rect 318586 280338 318822 280574
rect 318266 244658 318502 244894
rect 318586 244658 318822 244894
rect 318266 244338 318502 244574
rect 318586 244338 318822 244574
rect 318266 208658 318502 208894
rect 318586 208658 318822 208894
rect 318266 208338 318502 208574
rect 318586 208338 318822 208574
rect 318266 172658 318502 172894
rect 318586 172658 318822 172894
rect 318266 172338 318502 172574
rect 318586 172338 318822 172574
rect 318266 136658 318502 136894
rect 318586 136658 318822 136894
rect 318266 136338 318502 136574
rect 318586 136338 318822 136574
rect 318266 100658 318502 100894
rect 318586 100658 318822 100894
rect 318266 100338 318502 100574
rect 318586 100338 318822 100574
rect 318266 64658 318502 64894
rect 318586 64658 318822 64894
rect 318266 64338 318502 64574
rect 318586 64338 318822 64574
rect 318266 28658 318502 28894
rect 318586 28658 318822 28894
rect 318266 28338 318502 28574
rect 318586 28338 318822 28574
rect 320826 704602 321062 704838
rect 321146 704602 321382 704838
rect 320826 704282 321062 704518
rect 321146 704282 321382 704518
rect 320826 687218 321062 687454
rect 321146 687218 321382 687454
rect 320826 686898 321062 687134
rect 321146 686898 321382 687134
rect 320826 651218 321062 651454
rect 321146 651218 321382 651454
rect 320826 650898 321062 651134
rect 321146 650898 321382 651134
rect 320826 615218 321062 615454
rect 321146 615218 321382 615454
rect 320826 614898 321062 615134
rect 321146 614898 321382 615134
rect 320826 579218 321062 579454
rect 321146 579218 321382 579454
rect 320826 578898 321062 579134
rect 321146 578898 321382 579134
rect 320826 543218 321062 543454
rect 321146 543218 321382 543454
rect 320826 542898 321062 543134
rect 321146 542898 321382 543134
rect 320826 507218 321062 507454
rect 321146 507218 321382 507454
rect 320826 506898 321062 507134
rect 321146 506898 321382 507134
rect 320826 471218 321062 471454
rect 321146 471218 321382 471454
rect 320826 470898 321062 471134
rect 321146 470898 321382 471134
rect 320826 435218 321062 435454
rect 321146 435218 321382 435454
rect 320826 434898 321062 435134
rect 321146 434898 321382 435134
rect 320826 399218 321062 399454
rect 321146 399218 321382 399454
rect 320826 398898 321062 399134
rect 321146 398898 321382 399134
rect 320826 363218 321062 363454
rect 321146 363218 321382 363454
rect 320826 362898 321062 363134
rect 321146 362898 321382 363134
rect 320826 327218 321062 327454
rect 321146 327218 321382 327454
rect 320826 326898 321062 327134
rect 321146 326898 321382 327134
rect 320826 291218 321062 291454
rect 321146 291218 321382 291454
rect 320826 290898 321062 291134
rect 321146 290898 321382 291134
rect 320826 255218 321062 255454
rect 321146 255218 321382 255454
rect 320826 254898 321062 255134
rect 321146 254898 321382 255134
rect 320826 219218 321062 219454
rect 321146 219218 321382 219454
rect 320826 218898 321062 219134
rect 321146 218898 321382 219134
rect 320826 183218 321062 183454
rect 321146 183218 321382 183454
rect 320826 182898 321062 183134
rect 321146 182898 321382 183134
rect 320826 147218 321062 147454
rect 321146 147218 321382 147454
rect 320826 146898 321062 147134
rect 321146 146898 321382 147134
rect 320826 111218 321062 111454
rect 321146 111218 321382 111454
rect 320826 110898 321062 111134
rect 321146 110898 321382 111134
rect 320826 75218 321062 75454
rect 321146 75218 321382 75454
rect 320826 74898 321062 75134
rect 321146 74898 321382 75134
rect 320826 39218 321062 39454
rect 321146 39218 321382 39454
rect 320826 38898 321062 39134
rect 321146 38898 321382 39134
rect 320826 3218 321062 3454
rect 321146 3218 321382 3454
rect 320826 2898 321062 3134
rect 321146 2898 321382 3134
rect 320826 -582 321062 -346
rect 321146 -582 321382 -346
rect 320826 -902 321062 -666
rect 321146 -902 321382 -666
rect 331986 710362 332222 710598
rect 332306 710362 332542 710598
rect 331986 710042 332222 710278
rect 332306 710042 332542 710278
rect 328266 708442 328502 708678
rect 328586 708442 328822 708678
rect 328266 708122 328502 708358
rect 328586 708122 328822 708358
rect 321986 680378 322222 680614
rect 322306 680378 322542 680614
rect 321986 680058 322222 680294
rect 322306 680058 322542 680294
rect 321986 644378 322222 644614
rect 322306 644378 322542 644614
rect 321986 644058 322222 644294
rect 322306 644058 322542 644294
rect 321986 608378 322222 608614
rect 322306 608378 322542 608614
rect 321986 608058 322222 608294
rect 322306 608058 322542 608294
rect 321986 572378 322222 572614
rect 322306 572378 322542 572614
rect 321986 572058 322222 572294
rect 322306 572058 322542 572294
rect 321986 536378 322222 536614
rect 322306 536378 322542 536614
rect 321986 536058 322222 536294
rect 322306 536058 322542 536294
rect 321986 500378 322222 500614
rect 322306 500378 322542 500614
rect 321986 500058 322222 500294
rect 322306 500058 322542 500294
rect 321986 464378 322222 464614
rect 322306 464378 322542 464614
rect 321986 464058 322222 464294
rect 322306 464058 322542 464294
rect 321986 428378 322222 428614
rect 322306 428378 322542 428614
rect 321986 428058 322222 428294
rect 322306 428058 322542 428294
rect 321986 392378 322222 392614
rect 322306 392378 322542 392614
rect 321986 392058 322222 392294
rect 322306 392058 322542 392294
rect 321986 356378 322222 356614
rect 322306 356378 322542 356614
rect 321986 356058 322222 356294
rect 322306 356058 322542 356294
rect 321986 320378 322222 320614
rect 322306 320378 322542 320614
rect 321986 320058 322222 320294
rect 322306 320058 322542 320294
rect 321986 284378 322222 284614
rect 322306 284378 322542 284614
rect 321986 284058 322222 284294
rect 322306 284058 322542 284294
rect 321986 248378 322222 248614
rect 322306 248378 322542 248614
rect 321986 248058 322222 248294
rect 322306 248058 322542 248294
rect 321986 212378 322222 212614
rect 322306 212378 322542 212614
rect 321986 212058 322222 212294
rect 322306 212058 322542 212294
rect 321986 176378 322222 176614
rect 322306 176378 322542 176614
rect 321986 176058 322222 176294
rect 322306 176058 322542 176294
rect 321986 140378 322222 140614
rect 322306 140378 322542 140614
rect 321986 140058 322222 140294
rect 322306 140058 322542 140294
rect 321986 104378 322222 104614
rect 322306 104378 322542 104614
rect 321986 104058 322222 104294
rect 322306 104058 322542 104294
rect 321986 68378 322222 68614
rect 322306 68378 322542 68614
rect 321986 68058 322222 68294
rect 322306 68058 322542 68294
rect 321986 32378 322222 32614
rect 322306 32378 322542 32614
rect 321986 32058 322222 32294
rect 322306 32058 322542 32294
rect 318266 -5382 318502 -5146
rect 318586 -5382 318822 -5146
rect 318266 -5702 318502 -5466
rect 318586 -5702 318822 -5466
rect 311986 -6342 312222 -6106
rect 312306 -6342 312542 -6106
rect 311986 -6662 312222 -6426
rect 312306 -6662 312542 -6426
rect 324546 706522 324782 706758
rect 324866 706522 325102 706758
rect 324546 706202 324782 706438
rect 324866 706202 325102 706438
rect 324546 690938 324782 691174
rect 324866 690938 325102 691174
rect 324546 690618 324782 690854
rect 324866 690618 325102 690854
rect 324546 654938 324782 655174
rect 324866 654938 325102 655174
rect 324546 654618 324782 654854
rect 324866 654618 325102 654854
rect 324546 618938 324782 619174
rect 324866 618938 325102 619174
rect 324546 618618 324782 618854
rect 324866 618618 325102 618854
rect 324546 582938 324782 583174
rect 324866 582938 325102 583174
rect 324546 582618 324782 582854
rect 324866 582618 325102 582854
rect 324546 546938 324782 547174
rect 324866 546938 325102 547174
rect 324546 546618 324782 546854
rect 324866 546618 325102 546854
rect 324546 510938 324782 511174
rect 324866 510938 325102 511174
rect 324546 510618 324782 510854
rect 324866 510618 325102 510854
rect 324546 474938 324782 475174
rect 324866 474938 325102 475174
rect 324546 474618 324782 474854
rect 324866 474618 325102 474854
rect 324546 438938 324782 439174
rect 324866 438938 325102 439174
rect 324546 438618 324782 438854
rect 324866 438618 325102 438854
rect 324546 402938 324782 403174
rect 324866 402938 325102 403174
rect 324546 402618 324782 402854
rect 324866 402618 325102 402854
rect 324546 366938 324782 367174
rect 324866 366938 325102 367174
rect 324546 366618 324782 366854
rect 324866 366618 325102 366854
rect 324546 330938 324782 331174
rect 324866 330938 325102 331174
rect 324546 330618 324782 330854
rect 324866 330618 325102 330854
rect 324546 294938 324782 295174
rect 324866 294938 325102 295174
rect 324546 294618 324782 294854
rect 324866 294618 325102 294854
rect 324546 258938 324782 259174
rect 324866 258938 325102 259174
rect 324546 258618 324782 258854
rect 324866 258618 325102 258854
rect 324546 222938 324782 223174
rect 324866 222938 325102 223174
rect 324546 222618 324782 222854
rect 324866 222618 325102 222854
rect 324546 186938 324782 187174
rect 324866 186938 325102 187174
rect 324546 186618 324782 186854
rect 324866 186618 325102 186854
rect 324546 150938 324782 151174
rect 324866 150938 325102 151174
rect 324546 150618 324782 150854
rect 324866 150618 325102 150854
rect 324546 114938 324782 115174
rect 324866 114938 325102 115174
rect 324546 114618 324782 114854
rect 324866 114618 325102 114854
rect 324546 78938 324782 79174
rect 324866 78938 325102 79174
rect 324546 78618 324782 78854
rect 324866 78618 325102 78854
rect 324546 42938 324782 43174
rect 324866 42938 325102 43174
rect 324546 42618 324782 42854
rect 324866 42618 325102 42854
rect 324546 6938 324782 7174
rect 324866 6938 325102 7174
rect 324546 6618 324782 6854
rect 324866 6618 325102 6854
rect 324546 -2502 324782 -2266
rect 324866 -2502 325102 -2266
rect 324546 -2822 324782 -2586
rect 324866 -2822 325102 -2586
rect 328266 694658 328502 694894
rect 328586 694658 328822 694894
rect 328266 694338 328502 694574
rect 328586 694338 328822 694574
rect 328266 658658 328502 658894
rect 328586 658658 328822 658894
rect 328266 658338 328502 658574
rect 328586 658338 328822 658574
rect 328266 622658 328502 622894
rect 328586 622658 328822 622894
rect 328266 622338 328502 622574
rect 328586 622338 328822 622574
rect 328266 586658 328502 586894
rect 328586 586658 328822 586894
rect 328266 586338 328502 586574
rect 328586 586338 328822 586574
rect 328266 550658 328502 550894
rect 328586 550658 328822 550894
rect 328266 550338 328502 550574
rect 328586 550338 328822 550574
rect 328266 514658 328502 514894
rect 328586 514658 328822 514894
rect 328266 514338 328502 514574
rect 328586 514338 328822 514574
rect 328266 478658 328502 478894
rect 328586 478658 328822 478894
rect 328266 478338 328502 478574
rect 328586 478338 328822 478574
rect 328266 442658 328502 442894
rect 328586 442658 328822 442894
rect 328266 442338 328502 442574
rect 328586 442338 328822 442574
rect 328266 406658 328502 406894
rect 328586 406658 328822 406894
rect 328266 406338 328502 406574
rect 328586 406338 328822 406574
rect 328266 370658 328502 370894
rect 328586 370658 328822 370894
rect 328266 370338 328502 370574
rect 328586 370338 328822 370574
rect 328266 334658 328502 334894
rect 328586 334658 328822 334894
rect 328266 334338 328502 334574
rect 328586 334338 328822 334574
rect 328266 298658 328502 298894
rect 328586 298658 328822 298894
rect 328266 298338 328502 298574
rect 328586 298338 328822 298574
rect 328266 262658 328502 262894
rect 328586 262658 328822 262894
rect 328266 262338 328502 262574
rect 328586 262338 328822 262574
rect 328266 226658 328502 226894
rect 328586 226658 328822 226894
rect 328266 226338 328502 226574
rect 328586 226338 328822 226574
rect 328266 190658 328502 190894
rect 328586 190658 328822 190894
rect 328266 190338 328502 190574
rect 328586 190338 328822 190574
rect 328266 154658 328502 154894
rect 328586 154658 328822 154894
rect 328266 154338 328502 154574
rect 328586 154338 328822 154574
rect 328266 118658 328502 118894
rect 328586 118658 328822 118894
rect 328266 118338 328502 118574
rect 328586 118338 328822 118574
rect 328266 82658 328502 82894
rect 328586 82658 328822 82894
rect 328266 82338 328502 82574
rect 328586 82338 328822 82574
rect 328266 46658 328502 46894
rect 328586 46658 328822 46894
rect 328266 46338 328502 46574
rect 328586 46338 328822 46574
rect 328266 10658 328502 10894
rect 328586 10658 328822 10894
rect 328266 10338 328502 10574
rect 328586 10338 328822 10574
rect 330826 705562 331062 705798
rect 331146 705562 331382 705798
rect 330826 705242 331062 705478
rect 331146 705242 331382 705478
rect 330826 669218 331062 669454
rect 331146 669218 331382 669454
rect 330826 668898 331062 669134
rect 331146 668898 331382 669134
rect 330826 633218 331062 633454
rect 331146 633218 331382 633454
rect 330826 632898 331062 633134
rect 331146 632898 331382 633134
rect 330826 597218 331062 597454
rect 331146 597218 331382 597454
rect 330826 596898 331062 597134
rect 331146 596898 331382 597134
rect 330826 561218 331062 561454
rect 331146 561218 331382 561454
rect 330826 560898 331062 561134
rect 331146 560898 331382 561134
rect 330826 525218 331062 525454
rect 331146 525218 331382 525454
rect 330826 524898 331062 525134
rect 331146 524898 331382 525134
rect 330826 489218 331062 489454
rect 331146 489218 331382 489454
rect 330826 488898 331062 489134
rect 331146 488898 331382 489134
rect 330826 453218 331062 453454
rect 331146 453218 331382 453454
rect 330826 452898 331062 453134
rect 331146 452898 331382 453134
rect 330826 417218 331062 417454
rect 331146 417218 331382 417454
rect 330826 416898 331062 417134
rect 331146 416898 331382 417134
rect 330826 381218 331062 381454
rect 331146 381218 331382 381454
rect 330826 380898 331062 381134
rect 331146 380898 331382 381134
rect 330826 345218 331062 345454
rect 331146 345218 331382 345454
rect 330826 344898 331062 345134
rect 331146 344898 331382 345134
rect 330826 309218 331062 309454
rect 331146 309218 331382 309454
rect 330826 308898 331062 309134
rect 331146 308898 331382 309134
rect 330826 273218 331062 273454
rect 331146 273218 331382 273454
rect 330826 272898 331062 273134
rect 331146 272898 331382 273134
rect 330826 237218 331062 237454
rect 331146 237218 331382 237454
rect 330826 236898 331062 237134
rect 331146 236898 331382 237134
rect 330826 201218 331062 201454
rect 331146 201218 331382 201454
rect 330826 200898 331062 201134
rect 331146 200898 331382 201134
rect 330826 165218 331062 165454
rect 331146 165218 331382 165454
rect 330826 164898 331062 165134
rect 331146 164898 331382 165134
rect 330826 129218 331062 129454
rect 331146 129218 331382 129454
rect 330826 128898 331062 129134
rect 331146 128898 331382 129134
rect 330826 93218 331062 93454
rect 331146 93218 331382 93454
rect 330826 92898 331062 93134
rect 331146 92898 331382 93134
rect 330826 57218 331062 57454
rect 331146 57218 331382 57454
rect 330826 56898 331062 57134
rect 331146 56898 331382 57134
rect 330826 21218 331062 21454
rect 331146 21218 331382 21454
rect 330826 20898 331062 21134
rect 331146 20898 331382 21134
rect 330826 -1542 331062 -1306
rect 331146 -1542 331382 -1306
rect 330826 -1862 331062 -1626
rect 331146 -1862 331382 -1626
rect 341986 711322 342222 711558
rect 342306 711322 342542 711558
rect 341986 711002 342222 711238
rect 342306 711002 342542 711238
rect 338266 709402 338502 709638
rect 338586 709402 338822 709638
rect 338266 709082 338502 709318
rect 338586 709082 338822 709318
rect 331986 698378 332222 698614
rect 332306 698378 332542 698614
rect 331986 698058 332222 698294
rect 332306 698058 332542 698294
rect 331986 662378 332222 662614
rect 332306 662378 332542 662614
rect 331986 662058 332222 662294
rect 332306 662058 332542 662294
rect 331986 626378 332222 626614
rect 332306 626378 332542 626614
rect 331986 626058 332222 626294
rect 332306 626058 332542 626294
rect 331986 590378 332222 590614
rect 332306 590378 332542 590614
rect 331986 590058 332222 590294
rect 332306 590058 332542 590294
rect 331986 554378 332222 554614
rect 332306 554378 332542 554614
rect 331986 554058 332222 554294
rect 332306 554058 332542 554294
rect 331986 518378 332222 518614
rect 332306 518378 332542 518614
rect 331986 518058 332222 518294
rect 332306 518058 332542 518294
rect 331986 482378 332222 482614
rect 332306 482378 332542 482614
rect 331986 482058 332222 482294
rect 332306 482058 332542 482294
rect 331986 446378 332222 446614
rect 332306 446378 332542 446614
rect 331986 446058 332222 446294
rect 332306 446058 332542 446294
rect 331986 410378 332222 410614
rect 332306 410378 332542 410614
rect 331986 410058 332222 410294
rect 332306 410058 332542 410294
rect 331986 374378 332222 374614
rect 332306 374378 332542 374614
rect 331986 374058 332222 374294
rect 332306 374058 332542 374294
rect 331986 338378 332222 338614
rect 332306 338378 332542 338614
rect 331986 338058 332222 338294
rect 332306 338058 332542 338294
rect 331986 302378 332222 302614
rect 332306 302378 332542 302614
rect 331986 302058 332222 302294
rect 332306 302058 332542 302294
rect 331986 266378 332222 266614
rect 332306 266378 332542 266614
rect 331986 266058 332222 266294
rect 332306 266058 332542 266294
rect 331986 230378 332222 230614
rect 332306 230378 332542 230614
rect 331986 230058 332222 230294
rect 332306 230058 332542 230294
rect 331986 194378 332222 194614
rect 332306 194378 332542 194614
rect 331986 194058 332222 194294
rect 332306 194058 332542 194294
rect 331986 158378 332222 158614
rect 332306 158378 332542 158614
rect 331986 158058 332222 158294
rect 332306 158058 332542 158294
rect 331986 122378 332222 122614
rect 332306 122378 332542 122614
rect 331986 122058 332222 122294
rect 332306 122058 332542 122294
rect 331986 86378 332222 86614
rect 332306 86378 332542 86614
rect 331986 86058 332222 86294
rect 332306 86058 332542 86294
rect 331986 50378 332222 50614
rect 332306 50378 332542 50614
rect 331986 50058 332222 50294
rect 332306 50058 332542 50294
rect 331986 14378 332222 14614
rect 332306 14378 332542 14614
rect 331986 14058 332222 14294
rect 332306 14058 332542 14294
rect 328266 -4422 328502 -4186
rect 328586 -4422 328822 -4186
rect 328266 -4742 328502 -4506
rect 328586 -4742 328822 -4506
rect 321986 -7302 322222 -7066
rect 322306 -7302 322542 -7066
rect 321986 -7622 322222 -7386
rect 322306 -7622 322542 -7386
rect 334546 707482 334782 707718
rect 334866 707482 335102 707718
rect 334546 707162 334782 707398
rect 334866 707162 335102 707398
rect 334546 672938 334782 673174
rect 334866 672938 335102 673174
rect 334546 672618 334782 672854
rect 334866 672618 335102 672854
rect 334546 636938 334782 637174
rect 334866 636938 335102 637174
rect 334546 636618 334782 636854
rect 334866 636618 335102 636854
rect 334546 600938 334782 601174
rect 334866 600938 335102 601174
rect 334546 600618 334782 600854
rect 334866 600618 335102 600854
rect 334546 564938 334782 565174
rect 334866 564938 335102 565174
rect 334546 564618 334782 564854
rect 334866 564618 335102 564854
rect 334546 528938 334782 529174
rect 334866 528938 335102 529174
rect 334546 528618 334782 528854
rect 334866 528618 335102 528854
rect 334546 492938 334782 493174
rect 334866 492938 335102 493174
rect 334546 492618 334782 492854
rect 334866 492618 335102 492854
rect 334546 456938 334782 457174
rect 334866 456938 335102 457174
rect 334546 456618 334782 456854
rect 334866 456618 335102 456854
rect 334546 420938 334782 421174
rect 334866 420938 335102 421174
rect 334546 420618 334782 420854
rect 334866 420618 335102 420854
rect 334546 384938 334782 385174
rect 334866 384938 335102 385174
rect 334546 384618 334782 384854
rect 334866 384618 335102 384854
rect 334546 348938 334782 349174
rect 334866 348938 335102 349174
rect 334546 348618 334782 348854
rect 334866 348618 335102 348854
rect 334546 312938 334782 313174
rect 334866 312938 335102 313174
rect 334546 312618 334782 312854
rect 334866 312618 335102 312854
rect 334546 276938 334782 277174
rect 334866 276938 335102 277174
rect 334546 276618 334782 276854
rect 334866 276618 335102 276854
rect 334546 240938 334782 241174
rect 334866 240938 335102 241174
rect 334546 240618 334782 240854
rect 334866 240618 335102 240854
rect 334546 204938 334782 205174
rect 334866 204938 335102 205174
rect 334546 204618 334782 204854
rect 334866 204618 335102 204854
rect 334546 168938 334782 169174
rect 334866 168938 335102 169174
rect 334546 168618 334782 168854
rect 334866 168618 335102 168854
rect 334546 132938 334782 133174
rect 334866 132938 335102 133174
rect 334546 132618 334782 132854
rect 334866 132618 335102 132854
rect 334546 96938 334782 97174
rect 334866 96938 335102 97174
rect 334546 96618 334782 96854
rect 334866 96618 335102 96854
rect 334546 60938 334782 61174
rect 334866 60938 335102 61174
rect 334546 60618 334782 60854
rect 334866 60618 335102 60854
rect 334546 24938 334782 25174
rect 334866 24938 335102 25174
rect 334546 24618 334782 24854
rect 334866 24618 335102 24854
rect 334546 -3462 334782 -3226
rect 334866 -3462 335102 -3226
rect 334546 -3782 334782 -3546
rect 334866 -3782 335102 -3546
rect 338266 676658 338502 676894
rect 338586 676658 338822 676894
rect 338266 676338 338502 676574
rect 338586 676338 338822 676574
rect 338266 640658 338502 640894
rect 338586 640658 338822 640894
rect 338266 640338 338502 640574
rect 338586 640338 338822 640574
rect 338266 604658 338502 604894
rect 338586 604658 338822 604894
rect 338266 604338 338502 604574
rect 338586 604338 338822 604574
rect 338266 568658 338502 568894
rect 338586 568658 338822 568894
rect 338266 568338 338502 568574
rect 338586 568338 338822 568574
rect 338266 532658 338502 532894
rect 338586 532658 338822 532894
rect 338266 532338 338502 532574
rect 338586 532338 338822 532574
rect 338266 496658 338502 496894
rect 338586 496658 338822 496894
rect 338266 496338 338502 496574
rect 338586 496338 338822 496574
rect 338266 460658 338502 460894
rect 338586 460658 338822 460894
rect 338266 460338 338502 460574
rect 338586 460338 338822 460574
rect 338266 424658 338502 424894
rect 338586 424658 338822 424894
rect 338266 424338 338502 424574
rect 338586 424338 338822 424574
rect 338266 388658 338502 388894
rect 338586 388658 338822 388894
rect 338266 388338 338502 388574
rect 338586 388338 338822 388574
rect 338266 352658 338502 352894
rect 338586 352658 338822 352894
rect 338266 352338 338502 352574
rect 338586 352338 338822 352574
rect 338266 316658 338502 316894
rect 338586 316658 338822 316894
rect 338266 316338 338502 316574
rect 338586 316338 338822 316574
rect 338266 280658 338502 280894
rect 338586 280658 338822 280894
rect 338266 280338 338502 280574
rect 338586 280338 338822 280574
rect 338266 244658 338502 244894
rect 338586 244658 338822 244894
rect 338266 244338 338502 244574
rect 338586 244338 338822 244574
rect 338266 208658 338502 208894
rect 338586 208658 338822 208894
rect 338266 208338 338502 208574
rect 338586 208338 338822 208574
rect 338266 172658 338502 172894
rect 338586 172658 338822 172894
rect 338266 172338 338502 172574
rect 338586 172338 338822 172574
rect 338266 136658 338502 136894
rect 338586 136658 338822 136894
rect 338266 136338 338502 136574
rect 338586 136338 338822 136574
rect 338266 100658 338502 100894
rect 338586 100658 338822 100894
rect 338266 100338 338502 100574
rect 338586 100338 338822 100574
rect 338266 64658 338502 64894
rect 338586 64658 338822 64894
rect 338266 64338 338502 64574
rect 338586 64338 338822 64574
rect 338266 28658 338502 28894
rect 338586 28658 338822 28894
rect 338266 28338 338502 28574
rect 338586 28338 338822 28574
rect 340826 704602 341062 704838
rect 341146 704602 341382 704838
rect 340826 704282 341062 704518
rect 341146 704282 341382 704518
rect 340826 687218 341062 687454
rect 341146 687218 341382 687454
rect 340826 686898 341062 687134
rect 341146 686898 341382 687134
rect 340826 651218 341062 651454
rect 341146 651218 341382 651454
rect 340826 650898 341062 651134
rect 341146 650898 341382 651134
rect 340826 615218 341062 615454
rect 341146 615218 341382 615454
rect 340826 614898 341062 615134
rect 341146 614898 341382 615134
rect 340826 579218 341062 579454
rect 341146 579218 341382 579454
rect 340826 578898 341062 579134
rect 341146 578898 341382 579134
rect 340826 543218 341062 543454
rect 341146 543218 341382 543454
rect 340826 542898 341062 543134
rect 341146 542898 341382 543134
rect 340826 507218 341062 507454
rect 341146 507218 341382 507454
rect 340826 506898 341062 507134
rect 341146 506898 341382 507134
rect 340826 471218 341062 471454
rect 341146 471218 341382 471454
rect 340826 470898 341062 471134
rect 341146 470898 341382 471134
rect 340826 435218 341062 435454
rect 341146 435218 341382 435454
rect 340826 434898 341062 435134
rect 341146 434898 341382 435134
rect 340826 399218 341062 399454
rect 341146 399218 341382 399454
rect 340826 398898 341062 399134
rect 341146 398898 341382 399134
rect 340826 363218 341062 363454
rect 341146 363218 341382 363454
rect 340826 362898 341062 363134
rect 341146 362898 341382 363134
rect 340826 327218 341062 327454
rect 341146 327218 341382 327454
rect 340826 326898 341062 327134
rect 341146 326898 341382 327134
rect 340826 291218 341062 291454
rect 341146 291218 341382 291454
rect 340826 290898 341062 291134
rect 341146 290898 341382 291134
rect 340826 255218 341062 255454
rect 341146 255218 341382 255454
rect 340826 254898 341062 255134
rect 341146 254898 341382 255134
rect 340826 219218 341062 219454
rect 341146 219218 341382 219454
rect 340826 218898 341062 219134
rect 341146 218898 341382 219134
rect 340826 183218 341062 183454
rect 341146 183218 341382 183454
rect 340826 182898 341062 183134
rect 341146 182898 341382 183134
rect 340826 147218 341062 147454
rect 341146 147218 341382 147454
rect 340826 146898 341062 147134
rect 341146 146898 341382 147134
rect 340826 111218 341062 111454
rect 341146 111218 341382 111454
rect 340826 110898 341062 111134
rect 341146 110898 341382 111134
rect 340826 75218 341062 75454
rect 341146 75218 341382 75454
rect 340826 74898 341062 75134
rect 341146 74898 341382 75134
rect 340826 39218 341062 39454
rect 341146 39218 341382 39454
rect 340826 38898 341062 39134
rect 341146 38898 341382 39134
rect 340826 3218 341062 3454
rect 341146 3218 341382 3454
rect 340826 2898 341062 3134
rect 341146 2898 341382 3134
rect 340826 -582 341062 -346
rect 341146 -582 341382 -346
rect 340826 -902 341062 -666
rect 341146 -902 341382 -666
rect 351986 710362 352222 710598
rect 352306 710362 352542 710598
rect 351986 710042 352222 710278
rect 352306 710042 352542 710278
rect 348266 708442 348502 708678
rect 348586 708442 348822 708678
rect 348266 708122 348502 708358
rect 348586 708122 348822 708358
rect 341986 680378 342222 680614
rect 342306 680378 342542 680614
rect 341986 680058 342222 680294
rect 342306 680058 342542 680294
rect 341986 644378 342222 644614
rect 342306 644378 342542 644614
rect 341986 644058 342222 644294
rect 342306 644058 342542 644294
rect 341986 608378 342222 608614
rect 342306 608378 342542 608614
rect 341986 608058 342222 608294
rect 342306 608058 342542 608294
rect 341986 572378 342222 572614
rect 342306 572378 342542 572614
rect 341986 572058 342222 572294
rect 342306 572058 342542 572294
rect 341986 536378 342222 536614
rect 342306 536378 342542 536614
rect 341986 536058 342222 536294
rect 342306 536058 342542 536294
rect 341986 500378 342222 500614
rect 342306 500378 342542 500614
rect 341986 500058 342222 500294
rect 342306 500058 342542 500294
rect 341986 464378 342222 464614
rect 342306 464378 342542 464614
rect 341986 464058 342222 464294
rect 342306 464058 342542 464294
rect 341986 428378 342222 428614
rect 342306 428378 342542 428614
rect 341986 428058 342222 428294
rect 342306 428058 342542 428294
rect 341986 392378 342222 392614
rect 342306 392378 342542 392614
rect 341986 392058 342222 392294
rect 342306 392058 342542 392294
rect 341986 356378 342222 356614
rect 342306 356378 342542 356614
rect 341986 356058 342222 356294
rect 342306 356058 342542 356294
rect 341986 320378 342222 320614
rect 342306 320378 342542 320614
rect 341986 320058 342222 320294
rect 342306 320058 342542 320294
rect 341986 284378 342222 284614
rect 342306 284378 342542 284614
rect 341986 284058 342222 284294
rect 342306 284058 342542 284294
rect 341986 248378 342222 248614
rect 342306 248378 342542 248614
rect 341986 248058 342222 248294
rect 342306 248058 342542 248294
rect 341986 212378 342222 212614
rect 342306 212378 342542 212614
rect 341986 212058 342222 212294
rect 342306 212058 342542 212294
rect 341986 176378 342222 176614
rect 342306 176378 342542 176614
rect 341986 176058 342222 176294
rect 342306 176058 342542 176294
rect 341986 140378 342222 140614
rect 342306 140378 342542 140614
rect 341986 140058 342222 140294
rect 342306 140058 342542 140294
rect 341986 104378 342222 104614
rect 342306 104378 342542 104614
rect 341986 104058 342222 104294
rect 342306 104058 342542 104294
rect 341986 68378 342222 68614
rect 342306 68378 342542 68614
rect 341986 68058 342222 68294
rect 342306 68058 342542 68294
rect 341986 32378 342222 32614
rect 342306 32378 342542 32614
rect 341986 32058 342222 32294
rect 342306 32058 342542 32294
rect 338266 -5382 338502 -5146
rect 338586 -5382 338822 -5146
rect 338266 -5702 338502 -5466
rect 338586 -5702 338822 -5466
rect 331986 -6342 332222 -6106
rect 332306 -6342 332542 -6106
rect 331986 -6662 332222 -6426
rect 332306 -6662 332542 -6426
rect 344546 706522 344782 706758
rect 344866 706522 345102 706758
rect 344546 706202 344782 706438
rect 344866 706202 345102 706438
rect 344546 690938 344782 691174
rect 344866 690938 345102 691174
rect 344546 690618 344782 690854
rect 344866 690618 345102 690854
rect 344546 654938 344782 655174
rect 344866 654938 345102 655174
rect 344546 654618 344782 654854
rect 344866 654618 345102 654854
rect 344546 618938 344782 619174
rect 344866 618938 345102 619174
rect 344546 618618 344782 618854
rect 344866 618618 345102 618854
rect 344546 582938 344782 583174
rect 344866 582938 345102 583174
rect 344546 582618 344782 582854
rect 344866 582618 345102 582854
rect 344546 546938 344782 547174
rect 344866 546938 345102 547174
rect 344546 546618 344782 546854
rect 344866 546618 345102 546854
rect 344546 510938 344782 511174
rect 344866 510938 345102 511174
rect 344546 510618 344782 510854
rect 344866 510618 345102 510854
rect 344546 474938 344782 475174
rect 344866 474938 345102 475174
rect 344546 474618 344782 474854
rect 344866 474618 345102 474854
rect 344546 438938 344782 439174
rect 344866 438938 345102 439174
rect 344546 438618 344782 438854
rect 344866 438618 345102 438854
rect 344546 402938 344782 403174
rect 344866 402938 345102 403174
rect 344546 402618 344782 402854
rect 344866 402618 345102 402854
rect 344546 366938 344782 367174
rect 344866 366938 345102 367174
rect 344546 366618 344782 366854
rect 344866 366618 345102 366854
rect 344546 330938 344782 331174
rect 344866 330938 345102 331174
rect 344546 330618 344782 330854
rect 344866 330618 345102 330854
rect 344546 294938 344782 295174
rect 344866 294938 345102 295174
rect 344546 294618 344782 294854
rect 344866 294618 345102 294854
rect 344546 258938 344782 259174
rect 344866 258938 345102 259174
rect 344546 258618 344782 258854
rect 344866 258618 345102 258854
rect 344546 222938 344782 223174
rect 344866 222938 345102 223174
rect 344546 222618 344782 222854
rect 344866 222618 345102 222854
rect 344546 186938 344782 187174
rect 344866 186938 345102 187174
rect 344546 186618 344782 186854
rect 344866 186618 345102 186854
rect 344546 150938 344782 151174
rect 344866 150938 345102 151174
rect 344546 150618 344782 150854
rect 344866 150618 345102 150854
rect 344546 114938 344782 115174
rect 344866 114938 345102 115174
rect 344546 114618 344782 114854
rect 344866 114618 345102 114854
rect 344546 78938 344782 79174
rect 344866 78938 345102 79174
rect 344546 78618 344782 78854
rect 344866 78618 345102 78854
rect 344546 42938 344782 43174
rect 344866 42938 345102 43174
rect 344546 42618 344782 42854
rect 344866 42618 345102 42854
rect 344546 6938 344782 7174
rect 344866 6938 345102 7174
rect 344546 6618 344782 6854
rect 344866 6618 345102 6854
rect 344546 -2502 344782 -2266
rect 344866 -2502 345102 -2266
rect 344546 -2822 344782 -2586
rect 344866 -2822 345102 -2586
rect 348266 694658 348502 694894
rect 348586 694658 348822 694894
rect 348266 694338 348502 694574
rect 348586 694338 348822 694574
rect 348266 658658 348502 658894
rect 348586 658658 348822 658894
rect 348266 658338 348502 658574
rect 348586 658338 348822 658574
rect 348266 622658 348502 622894
rect 348586 622658 348822 622894
rect 348266 622338 348502 622574
rect 348586 622338 348822 622574
rect 348266 586658 348502 586894
rect 348586 586658 348822 586894
rect 348266 586338 348502 586574
rect 348586 586338 348822 586574
rect 348266 550658 348502 550894
rect 348586 550658 348822 550894
rect 348266 550338 348502 550574
rect 348586 550338 348822 550574
rect 348266 514658 348502 514894
rect 348586 514658 348822 514894
rect 348266 514338 348502 514574
rect 348586 514338 348822 514574
rect 348266 478658 348502 478894
rect 348586 478658 348822 478894
rect 348266 478338 348502 478574
rect 348586 478338 348822 478574
rect 348266 442658 348502 442894
rect 348586 442658 348822 442894
rect 348266 442338 348502 442574
rect 348586 442338 348822 442574
rect 348266 406658 348502 406894
rect 348586 406658 348822 406894
rect 348266 406338 348502 406574
rect 348586 406338 348822 406574
rect 348266 370658 348502 370894
rect 348586 370658 348822 370894
rect 348266 370338 348502 370574
rect 348586 370338 348822 370574
rect 348266 334658 348502 334894
rect 348586 334658 348822 334894
rect 348266 334338 348502 334574
rect 348586 334338 348822 334574
rect 348266 298658 348502 298894
rect 348586 298658 348822 298894
rect 348266 298338 348502 298574
rect 348586 298338 348822 298574
rect 348266 262658 348502 262894
rect 348586 262658 348822 262894
rect 348266 262338 348502 262574
rect 348586 262338 348822 262574
rect 348266 226658 348502 226894
rect 348586 226658 348822 226894
rect 348266 226338 348502 226574
rect 348586 226338 348822 226574
rect 348266 190658 348502 190894
rect 348586 190658 348822 190894
rect 348266 190338 348502 190574
rect 348586 190338 348822 190574
rect 348266 154658 348502 154894
rect 348586 154658 348822 154894
rect 348266 154338 348502 154574
rect 348586 154338 348822 154574
rect 348266 118658 348502 118894
rect 348586 118658 348822 118894
rect 348266 118338 348502 118574
rect 348586 118338 348822 118574
rect 348266 82658 348502 82894
rect 348586 82658 348822 82894
rect 348266 82338 348502 82574
rect 348586 82338 348822 82574
rect 348266 46658 348502 46894
rect 348586 46658 348822 46894
rect 348266 46338 348502 46574
rect 348586 46338 348822 46574
rect 348266 10658 348502 10894
rect 348586 10658 348822 10894
rect 348266 10338 348502 10574
rect 348586 10338 348822 10574
rect 350826 705562 351062 705798
rect 351146 705562 351382 705798
rect 350826 705242 351062 705478
rect 351146 705242 351382 705478
rect 350826 669218 351062 669454
rect 351146 669218 351382 669454
rect 350826 668898 351062 669134
rect 351146 668898 351382 669134
rect 350826 633218 351062 633454
rect 351146 633218 351382 633454
rect 350826 632898 351062 633134
rect 351146 632898 351382 633134
rect 350826 597218 351062 597454
rect 351146 597218 351382 597454
rect 350826 596898 351062 597134
rect 351146 596898 351382 597134
rect 350826 561218 351062 561454
rect 351146 561218 351382 561454
rect 350826 560898 351062 561134
rect 351146 560898 351382 561134
rect 350826 525218 351062 525454
rect 351146 525218 351382 525454
rect 350826 524898 351062 525134
rect 351146 524898 351382 525134
rect 350826 489218 351062 489454
rect 351146 489218 351382 489454
rect 350826 488898 351062 489134
rect 351146 488898 351382 489134
rect 350826 453218 351062 453454
rect 351146 453218 351382 453454
rect 350826 452898 351062 453134
rect 351146 452898 351382 453134
rect 350826 417218 351062 417454
rect 351146 417218 351382 417454
rect 350826 416898 351062 417134
rect 351146 416898 351382 417134
rect 350826 381218 351062 381454
rect 351146 381218 351382 381454
rect 350826 380898 351062 381134
rect 351146 380898 351382 381134
rect 350826 345218 351062 345454
rect 351146 345218 351382 345454
rect 350826 344898 351062 345134
rect 351146 344898 351382 345134
rect 350826 309218 351062 309454
rect 351146 309218 351382 309454
rect 350826 308898 351062 309134
rect 351146 308898 351382 309134
rect 350826 273218 351062 273454
rect 351146 273218 351382 273454
rect 350826 272898 351062 273134
rect 351146 272898 351382 273134
rect 350826 237218 351062 237454
rect 351146 237218 351382 237454
rect 350826 236898 351062 237134
rect 351146 236898 351382 237134
rect 350826 201218 351062 201454
rect 351146 201218 351382 201454
rect 350826 200898 351062 201134
rect 351146 200898 351382 201134
rect 350826 165218 351062 165454
rect 351146 165218 351382 165454
rect 350826 164898 351062 165134
rect 351146 164898 351382 165134
rect 350826 129218 351062 129454
rect 351146 129218 351382 129454
rect 350826 128898 351062 129134
rect 351146 128898 351382 129134
rect 350826 93218 351062 93454
rect 351146 93218 351382 93454
rect 350826 92898 351062 93134
rect 351146 92898 351382 93134
rect 350826 57218 351062 57454
rect 351146 57218 351382 57454
rect 350826 56898 351062 57134
rect 351146 56898 351382 57134
rect 350826 21218 351062 21454
rect 351146 21218 351382 21454
rect 350826 20898 351062 21134
rect 351146 20898 351382 21134
rect 350826 -1542 351062 -1306
rect 351146 -1542 351382 -1306
rect 350826 -1862 351062 -1626
rect 351146 -1862 351382 -1626
rect 361986 711322 362222 711558
rect 362306 711322 362542 711558
rect 361986 711002 362222 711238
rect 362306 711002 362542 711238
rect 358266 709402 358502 709638
rect 358586 709402 358822 709638
rect 358266 709082 358502 709318
rect 358586 709082 358822 709318
rect 351986 698378 352222 698614
rect 352306 698378 352542 698614
rect 351986 698058 352222 698294
rect 352306 698058 352542 698294
rect 351986 662378 352222 662614
rect 352306 662378 352542 662614
rect 351986 662058 352222 662294
rect 352306 662058 352542 662294
rect 351986 626378 352222 626614
rect 352306 626378 352542 626614
rect 351986 626058 352222 626294
rect 352306 626058 352542 626294
rect 351986 590378 352222 590614
rect 352306 590378 352542 590614
rect 351986 590058 352222 590294
rect 352306 590058 352542 590294
rect 351986 554378 352222 554614
rect 352306 554378 352542 554614
rect 351986 554058 352222 554294
rect 352306 554058 352542 554294
rect 351986 518378 352222 518614
rect 352306 518378 352542 518614
rect 351986 518058 352222 518294
rect 352306 518058 352542 518294
rect 351986 482378 352222 482614
rect 352306 482378 352542 482614
rect 351986 482058 352222 482294
rect 352306 482058 352542 482294
rect 351986 446378 352222 446614
rect 352306 446378 352542 446614
rect 351986 446058 352222 446294
rect 352306 446058 352542 446294
rect 351986 410378 352222 410614
rect 352306 410378 352542 410614
rect 351986 410058 352222 410294
rect 352306 410058 352542 410294
rect 351986 374378 352222 374614
rect 352306 374378 352542 374614
rect 351986 374058 352222 374294
rect 352306 374058 352542 374294
rect 351986 338378 352222 338614
rect 352306 338378 352542 338614
rect 351986 338058 352222 338294
rect 352306 338058 352542 338294
rect 351986 302378 352222 302614
rect 352306 302378 352542 302614
rect 351986 302058 352222 302294
rect 352306 302058 352542 302294
rect 351986 266378 352222 266614
rect 352306 266378 352542 266614
rect 351986 266058 352222 266294
rect 352306 266058 352542 266294
rect 351986 230378 352222 230614
rect 352306 230378 352542 230614
rect 351986 230058 352222 230294
rect 352306 230058 352542 230294
rect 351986 194378 352222 194614
rect 352306 194378 352542 194614
rect 351986 194058 352222 194294
rect 352306 194058 352542 194294
rect 351986 158378 352222 158614
rect 352306 158378 352542 158614
rect 351986 158058 352222 158294
rect 352306 158058 352542 158294
rect 351986 122378 352222 122614
rect 352306 122378 352542 122614
rect 351986 122058 352222 122294
rect 352306 122058 352542 122294
rect 351986 86378 352222 86614
rect 352306 86378 352542 86614
rect 351986 86058 352222 86294
rect 352306 86058 352542 86294
rect 351986 50378 352222 50614
rect 352306 50378 352542 50614
rect 351986 50058 352222 50294
rect 352306 50058 352542 50294
rect 351986 14378 352222 14614
rect 352306 14378 352542 14614
rect 351986 14058 352222 14294
rect 352306 14058 352542 14294
rect 348266 -4422 348502 -4186
rect 348586 -4422 348822 -4186
rect 348266 -4742 348502 -4506
rect 348586 -4742 348822 -4506
rect 341986 -7302 342222 -7066
rect 342306 -7302 342542 -7066
rect 341986 -7622 342222 -7386
rect 342306 -7622 342542 -7386
rect 354546 707482 354782 707718
rect 354866 707482 355102 707718
rect 354546 707162 354782 707398
rect 354866 707162 355102 707398
rect 354546 672938 354782 673174
rect 354866 672938 355102 673174
rect 354546 672618 354782 672854
rect 354866 672618 355102 672854
rect 354546 636938 354782 637174
rect 354866 636938 355102 637174
rect 354546 636618 354782 636854
rect 354866 636618 355102 636854
rect 354546 600938 354782 601174
rect 354866 600938 355102 601174
rect 354546 600618 354782 600854
rect 354866 600618 355102 600854
rect 354546 564938 354782 565174
rect 354866 564938 355102 565174
rect 354546 564618 354782 564854
rect 354866 564618 355102 564854
rect 354546 528938 354782 529174
rect 354866 528938 355102 529174
rect 354546 528618 354782 528854
rect 354866 528618 355102 528854
rect 354546 492938 354782 493174
rect 354866 492938 355102 493174
rect 354546 492618 354782 492854
rect 354866 492618 355102 492854
rect 354546 456938 354782 457174
rect 354866 456938 355102 457174
rect 354546 456618 354782 456854
rect 354866 456618 355102 456854
rect 354546 420938 354782 421174
rect 354866 420938 355102 421174
rect 354546 420618 354782 420854
rect 354866 420618 355102 420854
rect 354546 384938 354782 385174
rect 354866 384938 355102 385174
rect 354546 384618 354782 384854
rect 354866 384618 355102 384854
rect 354546 348938 354782 349174
rect 354866 348938 355102 349174
rect 354546 348618 354782 348854
rect 354866 348618 355102 348854
rect 354546 312938 354782 313174
rect 354866 312938 355102 313174
rect 354546 312618 354782 312854
rect 354866 312618 355102 312854
rect 354546 276938 354782 277174
rect 354866 276938 355102 277174
rect 354546 276618 354782 276854
rect 354866 276618 355102 276854
rect 354546 240938 354782 241174
rect 354866 240938 355102 241174
rect 354546 240618 354782 240854
rect 354866 240618 355102 240854
rect 354546 204938 354782 205174
rect 354866 204938 355102 205174
rect 354546 204618 354782 204854
rect 354866 204618 355102 204854
rect 354546 168938 354782 169174
rect 354866 168938 355102 169174
rect 354546 168618 354782 168854
rect 354866 168618 355102 168854
rect 354546 132938 354782 133174
rect 354866 132938 355102 133174
rect 354546 132618 354782 132854
rect 354866 132618 355102 132854
rect 354546 96938 354782 97174
rect 354866 96938 355102 97174
rect 354546 96618 354782 96854
rect 354866 96618 355102 96854
rect 354546 60938 354782 61174
rect 354866 60938 355102 61174
rect 354546 60618 354782 60854
rect 354866 60618 355102 60854
rect 354546 24938 354782 25174
rect 354866 24938 355102 25174
rect 354546 24618 354782 24854
rect 354866 24618 355102 24854
rect 354546 -3462 354782 -3226
rect 354866 -3462 355102 -3226
rect 354546 -3782 354782 -3546
rect 354866 -3782 355102 -3546
rect 358266 676658 358502 676894
rect 358586 676658 358822 676894
rect 358266 676338 358502 676574
rect 358586 676338 358822 676574
rect 358266 640658 358502 640894
rect 358586 640658 358822 640894
rect 358266 640338 358502 640574
rect 358586 640338 358822 640574
rect 358266 604658 358502 604894
rect 358586 604658 358822 604894
rect 358266 604338 358502 604574
rect 358586 604338 358822 604574
rect 358266 568658 358502 568894
rect 358586 568658 358822 568894
rect 358266 568338 358502 568574
rect 358586 568338 358822 568574
rect 358266 532658 358502 532894
rect 358586 532658 358822 532894
rect 358266 532338 358502 532574
rect 358586 532338 358822 532574
rect 358266 496658 358502 496894
rect 358586 496658 358822 496894
rect 358266 496338 358502 496574
rect 358586 496338 358822 496574
rect 358266 460658 358502 460894
rect 358586 460658 358822 460894
rect 358266 460338 358502 460574
rect 358586 460338 358822 460574
rect 358266 424658 358502 424894
rect 358586 424658 358822 424894
rect 358266 424338 358502 424574
rect 358586 424338 358822 424574
rect 358266 388658 358502 388894
rect 358586 388658 358822 388894
rect 358266 388338 358502 388574
rect 358586 388338 358822 388574
rect 358266 352658 358502 352894
rect 358586 352658 358822 352894
rect 358266 352338 358502 352574
rect 358586 352338 358822 352574
rect 358266 316658 358502 316894
rect 358586 316658 358822 316894
rect 358266 316338 358502 316574
rect 358586 316338 358822 316574
rect 358266 280658 358502 280894
rect 358586 280658 358822 280894
rect 358266 280338 358502 280574
rect 358586 280338 358822 280574
rect 358266 244658 358502 244894
rect 358586 244658 358822 244894
rect 358266 244338 358502 244574
rect 358586 244338 358822 244574
rect 358266 208658 358502 208894
rect 358586 208658 358822 208894
rect 358266 208338 358502 208574
rect 358586 208338 358822 208574
rect 358266 172658 358502 172894
rect 358586 172658 358822 172894
rect 358266 172338 358502 172574
rect 358586 172338 358822 172574
rect 358266 136658 358502 136894
rect 358586 136658 358822 136894
rect 358266 136338 358502 136574
rect 358586 136338 358822 136574
rect 358266 100658 358502 100894
rect 358586 100658 358822 100894
rect 358266 100338 358502 100574
rect 358586 100338 358822 100574
rect 358266 64658 358502 64894
rect 358586 64658 358822 64894
rect 358266 64338 358502 64574
rect 358586 64338 358822 64574
rect 358266 28658 358502 28894
rect 358586 28658 358822 28894
rect 358266 28338 358502 28574
rect 358586 28338 358822 28574
rect 360826 704602 361062 704838
rect 361146 704602 361382 704838
rect 360826 704282 361062 704518
rect 361146 704282 361382 704518
rect 360826 687218 361062 687454
rect 361146 687218 361382 687454
rect 360826 686898 361062 687134
rect 361146 686898 361382 687134
rect 360826 651218 361062 651454
rect 361146 651218 361382 651454
rect 360826 650898 361062 651134
rect 361146 650898 361382 651134
rect 360826 615218 361062 615454
rect 361146 615218 361382 615454
rect 360826 614898 361062 615134
rect 361146 614898 361382 615134
rect 360826 579218 361062 579454
rect 361146 579218 361382 579454
rect 360826 578898 361062 579134
rect 361146 578898 361382 579134
rect 360826 543218 361062 543454
rect 361146 543218 361382 543454
rect 360826 542898 361062 543134
rect 361146 542898 361382 543134
rect 360826 507218 361062 507454
rect 361146 507218 361382 507454
rect 360826 506898 361062 507134
rect 361146 506898 361382 507134
rect 360826 471218 361062 471454
rect 361146 471218 361382 471454
rect 360826 470898 361062 471134
rect 361146 470898 361382 471134
rect 360826 435218 361062 435454
rect 361146 435218 361382 435454
rect 360826 434898 361062 435134
rect 361146 434898 361382 435134
rect 360826 399218 361062 399454
rect 361146 399218 361382 399454
rect 360826 398898 361062 399134
rect 361146 398898 361382 399134
rect 360826 363218 361062 363454
rect 361146 363218 361382 363454
rect 360826 362898 361062 363134
rect 361146 362898 361382 363134
rect 360826 327218 361062 327454
rect 361146 327218 361382 327454
rect 360826 326898 361062 327134
rect 361146 326898 361382 327134
rect 360826 291218 361062 291454
rect 361146 291218 361382 291454
rect 360826 290898 361062 291134
rect 361146 290898 361382 291134
rect 360826 255218 361062 255454
rect 361146 255218 361382 255454
rect 360826 254898 361062 255134
rect 361146 254898 361382 255134
rect 360826 219218 361062 219454
rect 361146 219218 361382 219454
rect 360826 218898 361062 219134
rect 361146 218898 361382 219134
rect 360826 183218 361062 183454
rect 361146 183218 361382 183454
rect 360826 182898 361062 183134
rect 361146 182898 361382 183134
rect 360826 147218 361062 147454
rect 361146 147218 361382 147454
rect 360826 146898 361062 147134
rect 361146 146898 361382 147134
rect 360826 111218 361062 111454
rect 361146 111218 361382 111454
rect 360826 110898 361062 111134
rect 361146 110898 361382 111134
rect 360826 75218 361062 75454
rect 361146 75218 361382 75454
rect 360826 74898 361062 75134
rect 361146 74898 361382 75134
rect 360826 39218 361062 39454
rect 361146 39218 361382 39454
rect 360826 38898 361062 39134
rect 361146 38898 361382 39134
rect 360826 3218 361062 3454
rect 361146 3218 361382 3454
rect 360826 2898 361062 3134
rect 361146 2898 361382 3134
rect 360826 -582 361062 -346
rect 361146 -582 361382 -346
rect 360826 -902 361062 -666
rect 361146 -902 361382 -666
rect 371986 710362 372222 710598
rect 372306 710362 372542 710598
rect 371986 710042 372222 710278
rect 372306 710042 372542 710278
rect 368266 708442 368502 708678
rect 368586 708442 368822 708678
rect 368266 708122 368502 708358
rect 368586 708122 368822 708358
rect 361986 680378 362222 680614
rect 362306 680378 362542 680614
rect 361986 680058 362222 680294
rect 362306 680058 362542 680294
rect 361986 644378 362222 644614
rect 362306 644378 362542 644614
rect 361986 644058 362222 644294
rect 362306 644058 362542 644294
rect 361986 608378 362222 608614
rect 362306 608378 362542 608614
rect 361986 608058 362222 608294
rect 362306 608058 362542 608294
rect 361986 572378 362222 572614
rect 362306 572378 362542 572614
rect 361986 572058 362222 572294
rect 362306 572058 362542 572294
rect 361986 536378 362222 536614
rect 362306 536378 362542 536614
rect 361986 536058 362222 536294
rect 362306 536058 362542 536294
rect 361986 500378 362222 500614
rect 362306 500378 362542 500614
rect 361986 500058 362222 500294
rect 362306 500058 362542 500294
rect 361986 464378 362222 464614
rect 362306 464378 362542 464614
rect 361986 464058 362222 464294
rect 362306 464058 362542 464294
rect 361986 428378 362222 428614
rect 362306 428378 362542 428614
rect 361986 428058 362222 428294
rect 362306 428058 362542 428294
rect 361986 392378 362222 392614
rect 362306 392378 362542 392614
rect 361986 392058 362222 392294
rect 362306 392058 362542 392294
rect 361986 356378 362222 356614
rect 362306 356378 362542 356614
rect 361986 356058 362222 356294
rect 362306 356058 362542 356294
rect 361986 320378 362222 320614
rect 362306 320378 362542 320614
rect 361986 320058 362222 320294
rect 362306 320058 362542 320294
rect 361986 284378 362222 284614
rect 362306 284378 362542 284614
rect 361986 284058 362222 284294
rect 362306 284058 362542 284294
rect 361986 248378 362222 248614
rect 362306 248378 362542 248614
rect 361986 248058 362222 248294
rect 362306 248058 362542 248294
rect 361986 212378 362222 212614
rect 362306 212378 362542 212614
rect 361986 212058 362222 212294
rect 362306 212058 362542 212294
rect 361986 176378 362222 176614
rect 362306 176378 362542 176614
rect 361986 176058 362222 176294
rect 362306 176058 362542 176294
rect 361986 140378 362222 140614
rect 362306 140378 362542 140614
rect 361986 140058 362222 140294
rect 362306 140058 362542 140294
rect 361986 104378 362222 104614
rect 362306 104378 362542 104614
rect 361986 104058 362222 104294
rect 362306 104058 362542 104294
rect 361986 68378 362222 68614
rect 362306 68378 362542 68614
rect 361986 68058 362222 68294
rect 362306 68058 362542 68294
rect 361986 32378 362222 32614
rect 362306 32378 362542 32614
rect 361986 32058 362222 32294
rect 362306 32058 362542 32294
rect 358266 -5382 358502 -5146
rect 358586 -5382 358822 -5146
rect 358266 -5702 358502 -5466
rect 358586 -5702 358822 -5466
rect 351986 -6342 352222 -6106
rect 352306 -6342 352542 -6106
rect 351986 -6662 352222 -6426
rect 352306 -6662 352542 -6426
rect 364546 706522 364782 706758
rect 364866 706522 365102 706758
rect 364546 706202 364782 706438
rect 364866 706202 365102 706438
rect 364546 690938 364782 691174
rect 364866 690938 365102 691174
rect 364546 690618 364782 690854
rect 364866 690618 365102 690854
rect 364546 654938 364782 655174
rect 364866 654938 365102 655174
rect 364546 654618 364782 654854
rect 364866 654618 365102 654854
rect 364546 618938 364782 619174
rect 364866 618938 365102 619174
rect 364546 618618 364782 618854
rect 364866 618618 365102 618854
rect 364546 582938 364782 583174
rect 364866 582938 365102 583174
rect 364546 582618 364782 582854
rect 364866 582618 365102 582854
rect 364546 546938 364782 547174
rect 364866 546938 365102 547174
rect 364546 546618 364782 546854
rect 364866 546618 365102 546854
rect 364546 510938 364782 511174
rect 364866 510938 365102 511174
rect 364546 510618 364782 510854
rect 364866 510618 365102 510854
rect 364546 474938 364782 475174
rect 364866 474938 365102 475174
rect 364546 474618 364782 474854
rect 364866 474618 365102 474854
rect 364546 438938 364782 439174
rect 364866 438938 365102 439174
rect 364546 438618 364782 438854
rect 364866 438618 365102 438854
rect 364546 402938 364782 403174
rect 364866 402938 365102 403174
rect 364546 402618 364782 402854
rect 364866 402618 365102 402854
rect 364546 366938 364782 367174
rect 364866 366938 365102 367174
rect 364546 366618 364782 366854
rect 364866 366618 365102 366854
rect 364546 330938 364782 331174
rect 364866 330938 365102 331174
rect 364546 330618 364782 330854
rect 364866 330618 365102 330854
rect 364546 294938 364782 295174
rect 364866 294938 365102 295174
rect 364546 294618 364782 294854
rect 364866 294618 365102 294854
rect 364546 258938 364782 259174
rect 364866 258938 365102 259174
rect 364546 258618 364782 258854
rect 364866 258618 365102 258854
rect 364546 222938 364782 223174
rect 364866 222938 365102 223174
rect 364546 222618 364782 222854
rect 364866 222618 365102 222854
rect 364546 186938 364782 187174
rect 364866 186938 365102 187174
rect 364546 186618 364782 186854
rect 364866 186618 365102 186854
rect 364546 150938 364782 151174
rect 364866 150938 365102 151174
rect 364546 150618 364782 150854
rect 364866 150618 365102 150854
rect 364546 114938 364782 115174
rect 364866 114938 365102 115174
rect 364546 114618 364782 114854
rect 364866 114618 365102 114854
rect 364546 78938 364782 79174
rect 364866 78938 365102 79174
rect 364546 78618 364782 78854
rect 364866 78618 365102 78854
rect 364546 42938 364782 43174
rect 364866 42938 365102 43174
rect 364546 42618 364782 42854
rect 364866 42618 365102 42854
rect 364546 6938 364782 7174
rect 364866 6938 365102 7174
rect 364546 6618 364782 6854
rect 364866 6618 365102 6854
rect 364546 -2502 364782 -2266
rect 364866 -2502 365102 -2266
rect 364546 -2822 364782 -2586
rect 364866 -2822 365102 -2586
rect 368266 694658 368502 694894
rect 368586 694658 368822 694894
rect 368266 694338 368502 694574
rect 368586 694338 368822 694574
rect 368266 658658 368502 658894
rect 368586 658658 368822 658894
rect 368266 658338 368502 658574
rect 368586 658338 368822 658574
rect 368266 622658 368502 622894
rect 368586 622658 368822 622894
rect 368266 622338 368502 622574
rect 368586 622338 368822 622574
rect 368266 586658 368502 586894
rect 368586 586658 368822 586894
rect 368266 586338 368502 586574
rect 368586 586338 368822 586574
rect 368266 550658 368502 550894
rect 368586 550658 368822 550894
rect 368266 550338 368502 550574
rect 368586 550338 368822 550574
rect 368266 514658 368502 514894
rect 368586 514658 368822 514894
rect 368266 514338 368502 514574
rect 368586 514338 368822 514574
rect 368266 478658 368502 478894
rect 368586 478658 368822 478894
rect 368266 478338 368502 478574
rect 368586 478338 368822 478574
rect 368266 442658 368502 442894
rect 368586 442658 368822 442894
rect 368266 442338 368502 442574
rect 368586 442338 368822 442574
rect 368266 406658 368502 406894
rect 368586 406658 368822 406894
rect 368266 406338 368502 406574
rect 368586 406338 368822 406574
rect 368266 370658 368502 370894
rect 368586 370658 368822 370894
rect 368266 370338 368502 370574
rect 368586 370338 368822 370574
rect 368266 334658 368502 334894
rect 368586 334658 368822 334894
rect 368266 334338 368502 334574
rect 368586 334338 368822 334574
rect 368266 298658 368502 298894
rect 368586 298658 368822 298894
rect 368266 298338 368502 298574
rect 368586 298338 368822 298574
rect 368266 262658 368502 262894
rect 368586 262658 368822 262894
rect 368266 262338 368502 262574
rect 368586 262338 368822 262574
rect 368266 226658 368502 226894
rect 368586 226658 368822 226894
rect 368266 226338 368502 226574
rect 368586 226338 368822 226574
rect 368266 190658 368502 190894
rect 368586 190658 368822 190894
rect 368266 190338 368502 190574
rect 368586 190338 368822 190574
rect 368266 154658 368502 154894
rect 368586 154658 368822 154894
rect 368266 154338 368502 154574
rect 368586 154338 368822 154574
rect 368266 118658 368502 118894
rect 368586 118658 368822 118894
rect 368266 118338 368502 118574
rect 368586 118338 368822 118574
rect 368266 82658 368502 82894
rect 368586 82658 368822 82894
rect 368266 82338 368502 82574
rect 368586 82338 368822 82574
rect 368266 46658 368502 46894
rect 368586 46658 368822 46894
rect 368266 46338 368502 46574
rect 368586 46338 368822 46574
rect 368266 10658 368502 10894
rect 368586 10658 368822 10894
rect 368266 10338 368502 10574
rect 368586 10338 368822 10574
rect 370826 705562 371062 705798
rect 371146 705562 371382 705798
rect 370826 705242 371062 705478
rect 371146 705242 371382 705478
rect 370826 669218 371062 669454
rect 371146 669218 371382 669454
rect 370826 668898 371062 669134
rect 371146 668898 371382 669134
rect 370826 633218 371062 633454
rect 371146 633218 371382 633454
rect 370826 632898 371062 633134
rect 371146 632898 371382 633134
rect 370826 597218 371062 597454
rect 371146 597218 371382 597454
rect 370826 596898 371062 597134
rect 371146 596898 371382 597134
rect 370826 561218 371062 561454
rect 371146 561218 371382 561454
rect 370826 560898 371062 561134
rect 371146 560898 371382 561134
rect 370826 525218 371062 525454
rect 371146 525218 371382 525454
rect 370826 524898 371062 525134
rect 371146 524898 371382 525134
rect 370826 489218 371062 489454
rect 371146 489218 371382 489454
rect 370826 488898 371062 489134
rect 371146 488898 371382 489134
rect 370826 453218 371062 453454
rect 371146 453218 371382 453454
rect 370826 452898 371062 453134
rect 371146 452898 371382 453134
rect 370826 417218 371062 417454
rect 371146 417218 371382 417454
rect 370826 416898 371062 417134
rect 371146 416898 371382 417134
rect 370826 381218 371062 381454
rect 371146 381218 371382 381454
rect 370826 380898 371062 381134
rect 371146 380898 371382 381134
rect 370826 345218 371062 345454
rect 371146 345218 371382 345454
rect 370826 344898 371062 345134
rect 371146 344898 371382 345134
rect 370826 309218 371062 309454
rect 371146 309218 371382 309454
rect 370826 308898 371062 309134
rect 371146 308898 371382 309134
rect 370826 273218 371062 273454
rect 371146 273218 371382 273454
rect 370826 272898 371062 273134
rect 371146 272898 371382 273134
rect 370826 237218 371062 237454
rect 371146 237218 371382 237454
rect 370826 236898 371062 237134
rect 371146 236898 371382 237134
rect 370826 201218 371062 201454
rect 371146 201218 371382 201454
rect 370826 200898 371062 201134
rect 371146 200898 371382 201134
rect 370826 165218 371062 165454
rect 371146 165218 371382 165454
rect 370826 164898 371062 165134
rect 371146 164898 371382 165134
rect 370826 129218 371062 129454
rect 371146 129218 371382 129454
rect 370826 128898 371062 129134
rect 371146 128898 371382 129134
rect 370826 93218 371062 93454
rect 371146 93218 371382 93454
rect 370826 92898 371062 93134
rect 371146 92898 371382 93134
rect 370826 57218 371062 57454
rect 371146 57218 371382 57454
rect 370826 56898 371062 57134
rect 371146 56898 371382 57134
rect 370826 21218 371062 21454
rect 371146 21218 371382 21454
rect 370826 20898 371062 21134
rect 371146 20898 371382 21134
rect 370826 -1542 371062 -1306
rect 371146 -1542 371382 -1306
rect 370826 -1862 371062 -1626
rect 371146 -1862 371382 -1626
rect 381986 711322 382222 711558
rect 382306 711322 382542 711558
rect 381986 711002 382222 711238
rect 382306 711002 382542 711238
rect 378266 709402 378502 709638
rect 378586 709402 378822 709638
rect 378266 709082 378502 709318
rect 378586 709082 378822 709318
rect 371986 698378 372222 698614
rect 372306 698378 372542 698614
rect 371986 698058 372222 698294
rect 372306 698058 372542 698294
rect 371986 662378 372222 662614
rect 372306 662378 372542 662614
rect 371986 662058 372222 662294
rect 372306 662058 372542 662294
rect 371986 626378 372222 626614
rect 372306 626378 372542 626614
rect 371986 626058 372222 626294
rect 372306 626058 372542 626294
rect 371986 590378 372222 590614
rect 372306 590378 372542 590614
rect 371986 590058 372222 590294
rect 372306 590058 372542 590294
rect 371986 554378 372222 554614
rect 372306 554378 372542 554614
rect 371986 554058 372222 554294
rect 372306 554058 372542 554294
rect 371986 518378 372222 518614
rect 372306 518378 372542 518614
rect 371986 518058 372222 518294
rect 372306 518058 372542 518294
rect 371986 482378 372222 482614
rect 372306 482378 372542 482614
rect 371986 482058 372222 482294
rect 372306 482058 372542 482294
rect 371986 446378 372222 446614
rect 372306 446378 372542 446614
rect 371986 446058 372222 446294
rect 372306 446058 372542 446294
rect 371986 410378 372222 410614
rect 372306 410378 372542 410614
rect 371986 410058 372222 410294
rect 372306 410058 372542 410294
rect 371986 374378 372222 374614
rect 372306 374378 372542 374614
rect 371986 374058 372222 374294
rect 372306 374058 372542 374294
rect 371986 338378 372222 338614
rect 372306 338378 372542 338614
rect 371986 338058 372222 338294
rect 372306 338058 372542 338294
rect 371986 302378 372222 302614
rect 372306 302378 372542 302614
rect 371986 302058 372222 302294
rect 372306 302058 372542 302294
rect 371986 266378 372222 266614
rect 372306 266378 372542 266614
rect 371986 266058 372222 266294
rect 372306 266058 372542 266294
rect 371986 230378 372222 230614
rect 372306 230378 372542 230614
rect 371986 230058 372222 230294
rect 372306 230058 372542 230294
rect 371986 194378 372222 194614
rect 372306 194378 372542 194614
rect 371986 194058 372222 194294
rect 372306 194058 372542 194294
rect 371986 158378 372222 158614
rect 372306 158378 372542 158614
rect 371986 158058 372222 158294
rect 372306 158058 372542 158294
rect 371986 122378 372222 122614
rect 372306 122378 372542 122614
rect 371986 122058 372222 122294
rect 372306 122058 372542 122294
rect 371986 86378 372222 86614
rect 372306 86378 372542 86614
rect 371986 86058 372222 86294
rect 372306 86058 372542 86294
rect 371986 50378 372222 50614
rect 372306 50378 372542 50614
rect 371986 50058 372222 50294
rect 372306 50058 372542 50294
rect 371986 14378 372222 14614
rect 372306 14378 372542 14614
rect 371986 14058 372222 14294
rect 372306 14058 372542 14294
rect 368266 -4422 368502 -4186
rect 368586 -4422 368822 -4186
rect 368266 -4742 368502 -4506
rect 368586 -4742 368822 -4506
rect 361986 -7302 362222 -7066
rect 362306 -7302 362542 -7066
rect 361986 -7622 362222 -7386
rect 362306 -7622 362542 -7386
rect 374546 707482 374782 707718
rect 374866 707482 375102 707718
rect 374546 707162 374782 707398
rect 374866 707162 375102 707398
rect 374546 672938 374782 673174
rect 374866 672938 375102 673174
rect 374546 672618 374782 672854
rect 374866 672618 375102 672854
rect 374546 636938 374782 637174
rect 374866 636938 375102 637174
rect 374546 636618 374782 636854
rect 374866 636618 375102 636854
rect 374546 600938 374782 601174
rect 374866 600938 375102 601174
rect 374546 600618 374782 600854
rect 374866 600618 375102 600854
rect 374546 564938 374782 565174
rect 374866 564938 375102 565174
rect 374546 564618 374782 564854
rect 374866 564618 375102 564854
rect 374546 528938 374782 529174
rect 374866 528938 375102 529174
rect 374546 528618 374782 528854
rect 374866 528618 375102 528854
rect 374546 492938 374782 493174
rect 374866 492938 375102 493174
rect 374546 492618 374782 492854
rect 374866 492618 375102 492854
rect 374546 456938 374782 457174
rect 374866 456938 375102 457174
rect 374546 456618 374782 456854
rect 374866 456618 375102 456854
rect 374546 420938 374782 421174
rect 374866 420938 375102 421174
rect 374546 420618 374782 420854
rect 374866 420618 375102 420854
rect 374546 384938 374782 385174
rect 374866 384938 375102 385174
rect 374546 384618 374782 384854
rect 374866 384618 375102 384854
rect 374546 348938 374782 349174
rect 374866 348938 375102 349174
rect 374546 348618 374782 348854
rect 374866 348618 375102 348854
rect 374546 312938 374782 313174
rect 374866 312938 375102 313174
rect 374546 312618 374782 312854
rect 374866 312618 375102 312854
rect 374546 276938 374782 277174
rect 374866 276938 375102 277174
rect 374546 276618 374782 276854
rect 374866 276618 375102 276854
rect 374546 240938 374782 241174
rect 374866 240938 375102 241174
rect 374546 240618 374782 240854
rect 374866 240618 375102 240854
rect 374546 204938 374782 205174
rect 374866 204938 375102 205174
rect 374546 204618 374782 204854
rect 374866 204618 375102 204854
rect 374546 168938 374782 169174
rect 374866 168938 375102 169174
rect 374546 168618 374782 168854
rect 374866 168618 375102 168854
rect 374546 132938 374782 133174
rect 374866 132938 375102 133174
rect 374546 132618 374782 132854
rect 374866 132618 375102 132854
rect 374546 96938 374782 97174
rect 374866 96938 375102 97174
rect 374546 96618 374782 96854
rect 374866 96618 375102 96854
rect 374546 60938 374782 61174
rect 374866 60938 375102 61174
rect 374546 60618 374782 60854
rect 374866 60618 375102 60854
rect 374546 24938 374782 25174
rect 374866 24938 375102 25174
rect 374546 24618 374782 24854
rect 374866 24618 375102 24854
rect 374546 -3462 374782 -3226
rect 374866 -3462 375102 -3226
rect 374546 -3782 374782 -3546
rect 374866 -3782 375102 -3546
rect 378266 676658 378502 676894
rect 378586 676658 378822 676894
rect 378266 676338 378502 676574
rect 378586 676338 378822 676574
rect 378266 640658 378502 640894
rect 378586 640658 378822 640894
rect 378266 640338 378502 640574
rect 378586 640338 378822 640574
rect 378266 604658 378502 604894
rect 378586 604658 378822 604894
rect 378266 604338 378502 604574
rect 378586 604338 378822 604574
rect 378266 568658 378502 568894
rect 378586 568658 378822 568894
rect 378266 568338 378502 568574
rect 378586 568338 378822 568574
rect 378266 532658 378502 532894
rect 378586 532658 378822 532894
rect 378266 532338 378502 532574
rect 378586 532338 378822 532574
rect 378266 496658 378502 496894
rect 378586 496658 378822 496894
rect 378266 496338 378502 496574
rect 378586 496338 378822 496574
rect 378266 460658 378502 460894
rect 378586 460658 378822 460894
rect 378266 460338 378502 460574
rect 378586 460338 378822 460574
rect 378266 424658 378502 424894
rect 378586 424658 378822 424894
rect 378266 424338 378502 424574
rect 378586 424338 378822 424574
rect 378266 388658 378502 388894
rect 378586 388658 378822 388894
rect 378266 388338 378502 388574
rect 378586 388338 378822 388574
rect 378266 352658 378502 352894
rect 378586 352658 378822 352894
rect 378266 352338 378502 352574
rect 378586 352338 378822 352574
rect 378266 316658 378502 316894
rect 378586 316658 378822 316894
rect 378266 316338 378502 316574
rect 378586 316338 378822 316574
rect 378266 280658 378502 280894
rect 378586 280658 378822 280894
rect 378266 280338 378502 280574
rect 378586 280338 378822 280574
rect 378266 244658 378502 244894
rect 378586 244658 378822 244894
rect 378266 244338 378502 244574
rect 378586 244338 378822 244574
rect 378266 208658 378502 208894
rect 378586 208658 378822 208894
rect 378266 208338 378502 208574
rect 378586 208338 378822 208574
rect 378266 172658 378502 172894
rect 378586 172658 378822 172894
rect 378266 172338 378502 172574
rect 378586 172338 378822 172574
rect 378266 136658 378502 136894
rect 378586 136658 378822 136894
rect 378266 136338 378502 136574
rect 378586 136338 378822 136574
rect 378266 100658 378502 100894
rect 378586 100658 378822 100894
rect 378266 100338 378502 100574
rect 378586 100338 378822 100574
rect 378266 64658 378502 64894
rect 378586 64658 378822 64894
rect 378266 64338 378502 64574
rect 378586 64338 378822 64574
rect 378266 28658 378502 28894
rect 378586 28658 378822 28894
rect 378266 28338 378502 28574
rect 378586 28338 378822 28574
rect 380826 704602 381062 704838
rect 381146 704602 381382 704838
rect 380826 704282 381062 704518
rect 381146 704282 381382 704518
rect 380826 687218 381062 687454
rect 381146 687218 381382 687454
rect 380826 686898 381062 687134
rect 381146 686898 381382 687134
rect 380826 651218 381062 651454
rect 381146 651218 381382 651454
rect 380826 650898 381062 651134
rect 381146 650898 381382 651134
rect 380826 615218 381062 615454
rect 381146 615218 381382 615454
rect 380826 614898 381062 615134
rect 381146 614898 381382 615134
rect 380826 579218 381062 579454
rect 381146 579218 381382 579454
rect 380826 578898 381062 579134
rect 381146 578898 381382 579134
rect 380826 543218 381062 543454
rect 381146 543218 381382 543454
rect 380826 542898 381062 543134
rect 381146 542898 381382 543134
rect 380826 507218 381062 507454
rect 381146 507218 381382 507454
rect 380826 506898 381062 507134
rect 381146 506898 381382 507134
rect 380826 471218 381062 471454
rect 381146 471218 381382 471454
rect 380826 470898 381062 471134
rect 381146 470898 381382 471134
rect 380826 435218 381062 435454
rect 381146 435218 381382 435454
rect 380826 434898 381062 435134
rect 381146 434898 381382 435134
rect 380826 399218 381062 399454
rect 381146 399218 381382 399454
rect 380826 398898 381062 399134
rect 381146 398898 381382 399134
rect 380826 363218 381062 363454
rect 381146 363218 381382 363454
rect 380826 362898 381062 363134
rect 381146 362898 381382 363134
rect 380826 327218 381062 327454
rect 381146 327218 381382 327454
rect 380826 326898 381062 327134
rect 381146 326898 381382 327134
rect 380826 291218 381062 291454
rect 381146 291218 381382 291454
rect 380826 290898 381062 291134
rect 381146 290898 381382 291134
rect 380826 255218 381062 255454
rect 381146 255218 381382 255454
rect 380826 254898 381062 255134
rect 381146 254898 381382 255134
rect 380826 219218 381062 219454
rect 381146 219218 381382 219454
rect 380826 218898 381062 219134
rect 381146 218898 381382 219134
rect 380826 183218 381062 183454
rect 381146 183218 381382 183454
rect 380826 182898 381062 183134
rect 381146 182898 381382 183134
rect 380826 147218 381062 147454
rect 381146 147218 381382 147454
rect 380826 146898 381062 147134
rect 381146 146898 381382 147134
rect 380826 111218 381062 111454
rect 381146 111218 381382 111454
rect 380826 110898 381062 111134
rect 381146 110898 381382 111134
rect 380826 75218 381062 75454
rect 381146 75218 381382 75454
rect 380826 74898 381062 75134
rect 381146 74898 381382 75134
rect 380826 39218 381062 39454
rect 381146 39218 381382 39454
rect 380826 38898 381062 39134
rect 381146 38898 381382 39134
rect 380826 3218 381062 3454
rect 381146 3218 381382 3454
rect 380826 2898 381062 3134
rect 381146 2898 381382 3134
rect 380826 -582 381062 -346
rect 381146 -582 381382 -346
rect 380826 -902 381062 -666
rect 381146 -902 381382 -666
rect 391986 710362 392222 710598
rect 392306 710362 392542 710598
rect 391986 710042 392222 710278
rect 392306 710042 392542 710278
rect 388266 708442 388502 708678
rect 388586 708442 388822 708678
rect 388266 708122 388502 708358
rect 388586 708122 388822 708358
rect 381986 680378 382222 680614
rect 382306 680378 382542 680614
rect 381986 680058 382222 680294
rect 382306 680058 382542 680294
rect 381986 644378 382222 644614
rect 382306 644378 382542 644614
rect 381986 644058 382222 644294
rect 382306 644058 382542 644294
rect 381986 608378 382222 608614
rect 382306 608378 382542 608614
rect 381986 608058 382222 608294
rect 382306 608058 382542 608294
rect 381986 572378 382222 572614
rect 382306 572378 382542 572614
rect 381986 572058 382222 572294
rect 382306 572058 382542 572294
rect 381986 536378 382222 536614
rect 382306 536378 382542 536614
rect 381986 536058 382222 536294
rect 382306 536058 382542 536294
rect 381986 500378 382222 500614
rect 382306 500378 382542 500614
rect 381986 500058 382222 500294
rect 382306 500058 382542 500294
rect 381986 464378 382222 464614
rect 382306 464378 382542 464614
rect 381986 464058 382222 464294
rect 382306 464058 382542 464294
rect 381986 428378 382222 428614
rect 382306 428378 382542 428614
rect 381986 428058 382222 428294
rect 382306 428058 382542 428294
rect 381986 392378 382222 392614
rect 382306 392378 382542 392614
rect 381986 392058 382222 392294
rect 382306 392058 382542 392294
rect 381986 356378 382222 356614
rect 382306 356378 382542 356614
rect 381986 356058 382222 356294
rect 382306 356058 382542 356294
rect 381986 320378 382222 320614
rect 382306 320378 382542 320614
rect 381986 320058 382222 320294
rect 382306 320058 382542 320294
rect 381986 284378 382222 284614
rect 382306 284378 382542 284614
rect 381986 284058 382222 284294
rect 382306 284058 382542 284294
rect 381986 248378 382222 248614
rect 382306 248378 382542 248614
rect 381986 248058 382222 248294
rect 382306 248058 382542 248294
rect 381986 212378 382222 212614
rect 382306 212378 382542 212614
rect 381986 212058 382222 212294
rect 382306 212058 382542 212294
rect 381986 176378 382222 176614
rect 382306 176378 382542 176614
rect 381986 176058 382222 176294
rect 382306 176058 382542 176294
rect 381986 140378 382222 140614
rect 382306 140378 382542 140614
rect 381986 140058 382222 140294
rect 382306 140058 382542 140294
rect 381986 104378 382222 104614
rect 382306 104378 382542 104614
rect 381986 104058 382222 104294
rect 382306 104058 382542 104294
rect 381986 68378 382222 68614
rect 382306 68378 382542 68614
rect 381986 68058 382222 68294
rect 382306 68058 382542 68294
rect 381986 32378 382222 32614
rect 382306 32378 382542 32614
rect 381986 32058 382222 32294
rect 382306 32058 382542 32294
rect 378266 -5382 378502 -5146
rect 378586 -5382 378822 -5146
rect 378266 -5702 378502 -5466
rect 378586 -5702 378822 -5466
rect 371986 -6342 372222 -6106
rect 372306 -6342 372542 -6106
rect 371986 -6662 372222 -6426
rect 372306 -6662 372542 -6426
rect 384546 706522 384782 706758
rect 384866 706522 385102 706758
rect 384546 706202 384782 706438
rect 384866 706202 385102 706438
rect 384546 690938 384782 691174
rect 384866 690938 385102 691174
rect 384546 690618 384782 690854
rect 384866 690618 385102 690854
rect 384546 654938 384782 655174
rect 384866 654938 385102 655174
rect 384546 654618 384782 654854
rect 384866 654618 385102 654854
rect 384546 618938 384782 619174
rect 384866 618938 385102 619174
rect 384546 618618 384782 618854
rect 384866 618618 385102 618854
rect 384546 582938 384782 583174
rect 384866 582938 385102 583174
rect 384546 582618 384782 582854
rect 384866 582618 385102 582854
rect 384546 546938 384782 547174
rect 384866 546938 385102 547174
rect 384546 546618 384782 546854
rect 384866 546618 385102 546854
rect 384546 510938 384782 511174
rect 384866 510938 385102 511174
rect 384546 510618 384782 510854
rect 384866 510618 385102 510854
rect 384546 474938 384782 475174
rect 384866 474938 385102 475174
rect 384546 474618 384782 474854
rect 384866 474618 385102 474854
rect 384546 438938 384782 439174
rect 384866 438938 385102 439174
rect 384546 438618 384782 438854
rect 384866 438618 385102 438854
rect 384546 402938 384782 403174
rect 384866 402938 385102 403174
rect 384546 402618 384782 402854
rect 384866 402618 385102 402854
rect 384546 366938 384782 367174
rect 384866 366938 385102 367174
rect 384546 366618 384782 366854
rect 384866 366618 385102 366854
rect 384546 330938 384782 331174
rect 384866 330938 385102 331174
rect 384546 330618 384782 330854
rect 384866 330618 385102 330854
rect 384546 294938 384782 295174
rect 384866 294938 385102 295174
rect 384546 294618 384782 294854
rect 384866 294618 385102 294854
rect 384546 258938 384782 259174
rect 384866 258938 385102 259174
rect 384546 258618 384782 258854
rect 384866 258618 385102 258854
rect 384546 222938 384782 223174
rect 384866 222938 385102 223174
rect 384546 222618 384782 222854
rect 384866 222618 385102 222854
rect 384546 186938 384782 187174
rect 384866 186938 385102 187174
rect 384546 186618 384782 186854
rect 384866 186618 385102 186854
rect 384546 150938 384782 151174
rect 384866 150938 385102 151174
rect 384546 150618 384782 150854
rect 384866 150618 385102 150854
rect 384546 114938 384782 115174
rect 384866 114938 385102 115174
rect 384546 114618 384782 114854
rect 384866 114618 385102 114854
rect 384546 78938 384782 79174
rect 384866 78938 385102 79174
rect 384546 78618 384782 78854
rect 384866 78618 385102 78854
rect 384546 42938 384782 43174
rect 384866 42938 385102 43174
rect 384546 42618 384782 42854
rect 384866 42618 385102 42854
rect 384546 6938 384782 7174
rect 384866 6938 385102 7174
rect 384546 6618 384782 6854
rect 384866 6618 385102 6854
rect 384546 -2502 384782 -2266
rect 384866 -2502 385102 -2266
rect 384546 -2822 384782 -2586
rect 384866 -2822 385102 -2586
rect 388266 694658 388502 694894
rect 388586 694658 388822 694894
rect 388266 694338 388502 694574
rect 388586 694338 388822 694574
rect 388266 658658 388502 658894
rect 388586 658658 388822 658894
rect 388266 658338 388502 658574
rect 388586 658338 388822 658574
rect 388266 622658 388502 622894
rect 388586 622658 388822 622894
rect 388266 622338 388502 622574
rect 388586 622338 388822 622574
rect 388266 586658 388502 586894
rect 388586 586658 388822 586894
rect 388266 586338 388502 586574
rect 388586 586338 388822 586574
rect 388266 550658 388502 550894
rect 388586 550658 388822 550894
rect 388266 550338 388502 550574
rect 388586 550338 388822 550574
rect 388266 514658 388502 514894
rect 388586 514658 388822 514894
rect 388266 514338 388502 514574
rect 388586 514338 388822 514574
rect 388266 478658 388502 478894
rect 388586 478658 388822 478894
rect 388266 478338 388502 478574
rect 388586 478338 388822 478574
rect 388266 442658 388502 442894
rect 388586 442658 388822 442894
rect 388266 442338 388502 442574
rect 388586 442338 388822 442574
rect 388266 406658 388502 406894
rect 388586 406658 388822 406894
rect 388266 406338 388502 406574
rect 388586 406338 388822 406574
rect 388266 370658 388502 370894
rect 388586 370658 388822 370894
rect 388266 370338 388502 370574
rect 388586 370338 388822 370574
rect 388266 334658 388502 334894
rect 388586 334658 388822 334894
rect 388266 334338 388502 334574
rect 388586 334338 388822 334574
rect 388266 298658 388502 298894
rect 388586 298658 388822 298894
rect 388266 298338 388502 298574
rect 388586 298338 388822 298574
rect 388266 262658 388502 262894
rect 388586 262658 388822 262894
rect 388266 262338 388502 262574
rect 388586 262338 388822 262574
rect 388266 226658 388502 226894
rect 388586 226658 388822 226894
rect 388266 226338 388502 226574
rect 388586 226338 388822 226574
rect 388266 190658 388502 190894
rect 388586 190658 388822 190894
rect 388266 190338 388502 190574
rect 388586 190338 388822 190574
rect 388266 154658 388502 154894
rect 388586 154658 388822 154894
rect 388266 154338 388502 154574
rect 388586 154338 388822 154574
rect 388266 118658 388502 118894
rect 388586 118658 388822 118894
rect 388266 118338 388502 118574
rect 388586 118338 388822 118574
rect 388266 82658 388502 82894
rect 388586 82658 388822 82894
rect 388266 82338 388502 82574
rect 388586 82338 388822 82574
rect 388266 46658 388502 46894
rect 388586 46658 388822 46894
rect 388266 46338 388502 46574
rect 388586 46338 388822 46574
rect 388266 10658 388502 10894
rect 388586 10658 388822 10894
rect 388266 10338 388502 10574
rect 388586 10338 388822 10574
rect 390826 705562 391062 705798
rect 391146 705562 391382 705798
rect 390826 705242 391062 705478
rect 391146 705242 391382 705478
rect 390826 669218 391062 669454
rect 391146 669218 391382 669454
rect 390826 668898 391062 669134
rect 391146 668898 391382 669134
rect 390826 633218 391062 633454
rect 391146 633218 391382 633454
rect 390826 632898 391062 633134
rect 391146 632898 391382 633134
rect 390826 597218 391062 597454
rect 391146 597218 391382 597454
rect 390826 596898 391062 597134
rect 391146 596898 391382 597134
rect 390826 561218 391062 561454
rect 391146 561218 391382 561454
rect 390826 560898 391062 561134
rect 391146 560898 391382 561134
rect 390826 525218 391062 525454
rect 391146 525218 391382 525454
rect 390826 524898 391062 525134
rect 391146 524898 391382 525134
rect 390826 489218 391062 489454
rect 391146 489218 391382 489454
rect 390826 488898 391062 489134
rect 391146 488898 391382 489134
rect 390826 453218 391062 453454
rect 391146 453218 391382 453454
rect 390826 452898 391062 453134
rect 391146 452898 391382 453134
rect 390826 417218 391062 417454
rect 391146 417218 391382 417454
rect 390826 416898 391062 417134
rect 391146 416898 391382 417134
rect 390826 381218 391062 381454
rect 391146 381218 391382 381454
rect 390826 380898 391062 381134
rect 391146 380898 391382 381134
rect 390826 345218 391062 345454
rect 391146 345218 391382 345454
rect 390826 344898 391062 345134
rect 391146 344898 391382 345134
rect 390826 309218 391062 309454
rect 391146 309218 391382 309454
rect 390826 308898 391062 309134
rect 391146 308898 391382 309134
rect 390826 273218 391062 273454
rect 391146 273218 391382 273454
rect 390826 272898 391062 273134
rect 391146 272898 391382 273134
rect 390826 237218 391062 237454
rect 391146 237218 391382 237454
rect 390826 236898 391062 237134
rect 391146 236898 391382 237134
rect 390826 201218 391062 201454
rect 391146 201218 391382 201454
rect 390826 200898 391062 201134
rect 391146 200898 391382 201134
rect 390826 165218 391062 165454
rect 391146 165218 391382 165454
rect 390826 164898 391062 165134
rect 391146 164898 391382 165134
rect 390826 129218 391062 129454
rect 391146 129218 391382 129454
rect 390826 128898 391062 129134
rect 391146 128898 391382 129134
rect 390826 93218 391062 93454
rect 391146 93218 391382 93454
rect 390826 92898 391062 93134
rect 391146 92898 391382 93134
rect 390826 57218 391062 57454
rect 391146 57218 391382 57454
rect 390826 56898 391062 57134
rect 391146 56898 391382 57134
rect 390826 21218 391062 21454
rect 391146 21218 391382 21454
rect 390826 20898 391062 21134
rect 391146 20898 391382 21134
rect 390826 -1542 391062 -1306
rect 391146 -1542 391382 -1306
rect 390826 -1862 391062 -1626
rect 391146 -1862 391382 -1626
rect 401986 711322 402222 711558
rect 402306 711322 402542 711558
rect 401986 711002 402222 711238
rect 402306 711002 402542 711238
rect 398266 709402 398502 709638
rect 398586 709402 398822 709638
rect 398266 709082 398502 709318
rect 398586 709082 398822 709318
rect 391986 698378 392222 698614
rect 392306 698378 392542 698614
rect 391986 698058 392222 698294
rect 392306 698058 392542 698294
rect 391986 662378 392222 662614
rect 392306 662378 392542 662614
rect 391986 662058 392222 662294
rect 392306 662058 392542 662294
rect 391986 626378 392222 626614
rect 392306 626378 392542 626614
rect 391986 626058 392222 626294
rect 392306 626058 392542 626294
rect 391986 590378 392222 590614
rect 392306 590378 392542 590614
rect 391986 590058 392222 590294
rect 392306 590058 392542 590294
rect 391986 554378 392222 554614
rect 392306 554378 392542 554614
rect 391986 554058 392222 554294
rect 392306 554058 392542 554294
rect 391986 518378 392222 518614
rect 392306 518378 392542 518614
rect 391986 518058 392222 518294
rect 392306 518058 392542 518294
rect 391986 482378 392222 482614
rect 392306 482378 392542 482614
rect 391986 482058 392222 482294
rect 392306 482058 392542 482294
rect 391986 446378 392222 446614
rect 392306 446378 392542 446614
rect 391986 446058 392222 446294
rect 392306 446058 392542 446294
rect 391986 410378 392222 410614
rect 392306 410378 392542 410614
rect 391986 410058 392222 410294
rect 392306 410058 392542 410294
rect 391986 374378 392222 374614
rect 392306 374378 392542 374614
rect 391986 374058 392222 374294
rect 392306 374058 392542 374294
rect 391986 338378 392222 338614
rect 392306 338378 392542 338614
rect 391986 338058 392222 338294
rect 392306 338058 392542 338294
rect 391986 302378 392222 302614
rect 392306 302378 392542 302614
rect 391986 302058 392222 302294
rect 392306 302058 392542 302294
rect 391986 266378 392222 266614
rect 392306 266378 392542 266614
rect 391986 266058 392222 266294
rect 392306 266058 392542 266294
rect 391986 230378 392222 230614
rect 392306 230378 392542 230614
rect 391986 230058 392222 230294
rect 392306 230058 392542 230294
rect 391986 194378 392222 194614
rect 392306 194378 392542 194614
rect 391986 194058 392222 194294
rect 392306 194058 392542 194294
rect 391986 158378 392222 158614
rect 392306 158378 392542 158614
rect 391986 158058 392222 158294
rect 392306 158058 392542 158294
rect 391986 122378 392222 122614
rect 392306 122378 392542 122614
rect 391986 122058 392222 122294
rect 392306 122058 392542 122294
rect 391986 86378 392222 86614
rect 392306 86378 392542 86614
rect 391986 86058 392222 86294
rect 392306 86058 392542 86294
rect 391986 50378 392222 50614
rect 392306 50378 392542 50614
rect 391986 50058 392222 50294
rect 392306 50058 392542 50294
rect 391986 14378 392222 14614
rect 392306 14378 392542 14614
rect 391986 14058 392222 14294
rect 392306 14058 392542 14294
rect 388266 -4422 388502 -4186
rect 388586 -4422 388822 -4186
rect 388266 -4742 388502 -4506
rect 388586 -4742 388822 -4506
rect 381986 -7302 382222 -7066
rect 382306 -7302 382542 -7066
rect 381986 -7622 382222 -7386
rect 382306 -7622 382542 -7386
rect 394546 707482 394782 707718
rect 394866 707482 395102 707718
rect 394546 707162 394782 707398
rect 394866 707162 395102 707398
rect 394546 672938 394782 673174
rect 394866 672938 395102 673174
rect 394546 672618 394782 672854
rect 394866 672618 395102 672854
rect 394546 636938 394782 637174
rect 394866 636938 395102 637174
rect 394546 636618 394782 636854
rect 394866 636618 395102 636854
rect 394546 600938 394782 601174
rect 394866 600938 395102 601174
rect 394546 600618 394782 600854
rect 394866 600618 395102 600854
rect 394546 564938 394782 565174
rect 394866 564938 395102 565174
rect 394546 564618 394782 564854
rect 394866 564618 395102 564854
rect 394546 528938 394782 529174
rect 394866 528938 395102 529174
rect 394546 528618 394782 528854
rect 394866 528618 395102 528854
rect 394546 492938 394782 493174
rect 394866 492938 395102 493174
rect 394546 492618 394782 492854
rect 394866 492618 395102 492854
rect 394546 456938 394782 457174
rect 394866 456938 395102 457174
rect 394546 456618 394782 456854
rect 394866 456618 395102 456854
rect 394546 420938 394782 421174
rect 394866 420938 395102 421174
rect 394546 420618 394782 420854
rect 394866 420618 395102 420854
rect 394546 384938 394782 385174
rect 394866 384938 395102 385174
rect 394546 384618 394782 384854
rect 394866 384618 395102 384854
rect 394546 348938 394782 349174
rect 394866 348938 395102 349174
rect 394546 348618 394782 348854
rect 394866 348618 395102 348854
rect 394546 312938 394782 313174
rect 394866 312938 395102 313174
rect 394546 312618 394782 312854
rect 394866 312618 395102 312854
rect 394546 276938 394782 277174
rect 394866 276938 395102 277174
rect 394546 276618 394782 276854
rect 394866 276618 395102 276854
rect 394546 240938 394782 241174
rect 394866 240938 395102 241174
rect 394546 240618 394782 240854
rect 394866 240618 395102 240854
rect 394546 204938 394782 205174
rect 394866 204938 395102 205174
rect 394546 204618 394782 204854
rect 394866 204618 395102 204854
rect 394546 168938 394782 169174
rect 394866 168938 395102 169174
rect 394546 168618 394782 168854
rect 394866 168618 395102 168854
rect 394546 132938 394782 133174
rect 394866 132938 395102 133174
rect 394546 132618 394782 132854
rect 394866 132618 395102 132854
rect 394546 96938 394782 97174
rect 394866 96938 395102 97174
rect 394546 96618 394782 96854
rect 394866 96618 395102 96854
rect 394546 60938 394782 61174
rect 394866 60938 395102 61174
rect 394546 60618 394782 60854
rect 394866 60618 395102 60854
rect 394546 24938 394782 25174
rect 394866 24938 395102 25174
rect 394546 24618 394782 24854
rect 394866 24618 395102 24854
rect 394546 -3462 394782 -3226
rect 394866 -3462 395102 -3226
rect 394546 -3782 394782 -3546
rect 394866 -3782 395102 -3546
rect 398266 676658 398502 676894
rect 398586 676658 398822 676894
rect 398266 676338 398502 676574
rect 398586 676338 398822 676574
rect 398266 640658 398502 640894
rect 398586 640658 398822 640894
rect 398266 640338 398502 640574
rect 398586 640338 398822 640574
rect 398266 604658 398502 604894
rect 398586 604658 398822 604894
rect 398266 604338 398502 604574
rect 398586 604338 398822 604574
rect 398266 568658 398502 568894
rect 398586 568658 398822 568894
rect 398266 568338 398502 568574
rect 398586 568338 398822 568574
rect 398266 532658 398502 532894
rect 398586 532658 398822 532894
rect 398266 532338 398502 532574
rect 398586 532338 398822 532574
rect 398266 496658 398502 496894
rect 398586 496658 398822 496894
rect 398266 496338 398502 496574
rect 398586 496338 398822 496574
rect 398266 460658 398502 460894
rect 398586 460658 398822 460894
rect 398266 460338 398502 460574
rect 398586 460338 398822 460574
rect 398266 424658 398502 424894
rect 398586 424658 398822 424894
rect 398266 424338 398502 424574
rect 398586 424338 398822 424574
rect 398266 388658 398502 388894
rect 398586 388658 398822 388894
rect 398266 388338 398502 388574
rect 398586 388338 398822 388574
rect 398266 352658 398502 352894
rect 398586 352658 398822 352894
rect 398266 352338 398502 352574
rect 398586 352338 398822 352574
rect 398266 316658 398502 316894
rect 398586 316658 398822 316894
rect 398266 316338 398502 316574
rect 398586 316338 398822 316574
rect 398266 280658 398502 280894
rect 398586 280658 398822 280894
rect 398266 280338 398502 280574
rect 398586 280338 398822 280574
rect 398266 244658 398502 244894
rect 398586 244658 398822 244894
rect 398266 244338 398502 244574
rect 398586 244338 398822 244574
rect 398266 208658 398502 208894
rect 398586 208658 398822 208894
rect 398266 208338 398502 208574
rect 398586 208338 398822 208574
rect 398266 172658 398502 172894
rect 398586 172658 398822 172894
rect 398266 172338 398502 172574
rect 398586 172338 398822 172574
rect 398266 136658 398502 136894
rect 398586 136658 398822 136894
rect 398266 136338 398502 136574
rect 398586 136338 398822 136574
rect 398266 100658 398502 100894
rect 398586 100658 398822 100894
rect 398266 100338 398502 100574
rect 398586 100338 398822 100574
rect 398266 64658 398502 64894
rect 398586 64658 398822 64894
rect 398266 64338 398502 64574
rect 398586 64338 398822 64574
rect 398266 28658 398502 28894
rect 398586 28658 398822 28894
rect 398266 28338 398502 28574
rect 398586 28338 398822 28574
rect 400826 704602 401062 704838
rect 401146 704602 401382 704838
rect 400826 704282 401062 704518
rect 401146 704282 401382 704518
rect 400826 687218 401062 687454
rect 401146 687218 401382 687454
rect 400826 686898 401062 687134
rect 401146 686898 401382 687134
rect 400826 651218 401062 651454
rect 401146 651218 401382 651454
rect 400826 650898 401062 651134
rect 401146 650898 401382 651134
rect 400826 615218 401062 615454
rect 401146 615218 401382 615454
rect 400826 614898 401062 615134
rect 401146 614898 401382 615134
rect 400826 579218 401062 579454
rect 401146 579218 401382 579454
rect 400826 578898 401062 579134
rect 401146 578898 401382 579134
rect 400826 543218 401062 543454
rect 401146 543218 401382 543454
rect 400826 542898 401062 543134
rect 401146 542898 401382 543134
rect 400826 507218 401062 507454
rect 401146 507218 401382 507454
rect 400826 506898 401062 507134
rect 401146 506898 401382 507134
rect 400826 471218 401062 471454
rect 401146 471218 401382 471454
rect 400826 470898 401062 471134
rect 401146 470898 401382 471134
rect 400826 435218 401062 435454
rect 401146 435218 401382 435454
rect 400826 434898 401062 435134
rect 401146 434898 401382 435134
rect 400826 399218 401062 399454
rect 401146 399218 401382 399454
rect 400826 398898 401062 399134
rect 401146 398898 401382 399134
rect 400826 363218 401062 363454
rect 401146 363218 401382 363454
rect 400826 362898 401062 363134
rect 401146 362898 401382 363134
rect 400826 327218 401062 327454
rect 401146 327218 401382 327454
rect 400826 326898 401062 327134
rect 401146 326898 401382 327134
rect 400826 291218 401062 291454
rect 401146 291218 401382 291454
rect 400826 290898 401062 291134
rect 401146 290898 401382 291134
rect 400826 255218 401062 255454
rect 401146 255218 401382 255454
rect 400826 254898 401062 255134
rect 401146 254898 401382 255134
rect 400826 219218 401062 219454
rect 401146 219218 401382 219454
rect 400826 218898 401062 219134
rect 401146 218898 401382 219134
rect 400826 183218 401062 183454
rect 401146 183218 401382 183454
rect 400826 182898 401062 183134
rect 401146 182898 401382 183134
rect 400826 147218 401062 147454
rect 401146 147218 401382 147454
rect 400826 146898 401062 147134
rect 401146 146898 401382 147134
rect 400826 111218 401062 111454
rect 401146 111218 401382 111454
rect 400826 110898 401062 111134
rect 401146 110898 401382 111134
rect 400826 75218 401062 75454
rect 401146 75218 401382 75454
rect 400826 74898 401062 75134
rect 401146 74898 401382 75134
rect 400826 39218 401062 39454
rect 401146 39218 401382 39454
rect 400826 38898 401062 39134
rect 401146 38898 401382 39134
rect 400826 3218 401062 3454
rect 401146 3218 401382 3454
rect 400826 2898 401062 3134
rect 401146 2898 401382 3134
rect 400826 -582 401062 -346
rect 401146 -582 401382 -346
rect 400826 -902 401062 -666
rect 401146 -902 401382 -666
rect 411986 710362 412222 710598
rect 412306 710362 412542 710598
rect 411986 710042 412222 710278
rect 412306 710042 412542 710278
rect 408266 708442 408502 708678
rect 408586 708442 408822 708678
rect 408266 708122 408502 708358
rect 408586 708122 408822 708358
rect 401986 680378 402222 680614
rect 402306 680378 402542 680614
rect 401986 680058 402222 680294
rect 402306 680058 402542 680294
rect 401986 644378 402222 644614
rect 402306 644378 402542 644614
rect 401986 644058 402222 644294
rect 402306 644058 402542 644294
rect 401986 608378 402222 608614
rect 402306 608378 402542 608614
rect 401986 608058 402222 608294
rect 402306 608058 402542 608294
rect 401986 572378 402222 572614
rect 402306 572378 402542 572614
rect 401986 572058 402222 572294
rect 402306 572058 402542 572294
rect 401986 536378 402222 536614
rect 402306 536378 402542 536614
rect 401986 536058 402222 536294
rect 402306 536058 402542 536294
rect 401986 500378 402222 500614
rect 402306 500378 402542 500614
rect 401986 500058 402222 500294
rect 402306 500058 402542 500294
rect 401986 464378 402222 464614
rect 402306 464378 402542 464614
rect 401986 464058 402222 464294
rect 402306 464058 402542 464294
rect 401986 428378 402222 428614
rect 402306 428378 402542 428614
rect 401986 428058 402222 428294
rect 402306 428058 402542 428294
rect 401986 392378 402222 392614
rect 402306 392378 402542 392614
rect 401986 392058 402222 392294
rect 402306 392058 402542 392294
rect 401986 356378 402222 356614
rect 402306 356378 402542 356614
rect 401986 356058 402222 356294
rect 402306 356058 402542 356294
rect 401986 320378 402222 320614
rect 402306 320378 402542 320614
rect 401986 320058 402222 320294
rect 402306 320058 402542 320294
rect 401986 284378 402222 284614
rect 402306 284378 402542 284614
rect 401986 284058 402222 284294
rect 402306 284058 402542 284294
rect 401986 248378 402222 248614
rect 402306 248378 402542 248614
rect 401986 248058 402222 248294
rect 402306 248058 402542 248294
rect 401986 212378 402222 212614
rect 402306 212378 402542 212614
rect 401986 212058 402222 212294
rect 402306 212058 402542 212294
rect 401986 176378 402222 176614
rect 402306 176378 402542 176614
rect 401986 176058 402222 176294
rect 402306 176058 402542 176294
rect 401986 140378 402222 140614
rect 402306 140378 402542 140614
rect 401986 140058 402222 140294
rect 402306 140058 402542 140294
rect 401986 104378 402222 104614
rect 402306 104378 402542 104614
rect 401986 104058 402222 104294
rect 402306 104058 402542 104294
rect 401986 68378 402222 68614
rect 402306 68378 402542 68614
rect 401986 68058 402222 68294
rect 402306 68058 402542 68294
rect 401986 32378 402222 32614
rect 402306 32378 402542 32614
rect 401986 32058 402222 32294
rect 402306 32058 402542 32294
rect 398266 -5382 398502 -5146
rect 398586 -5382 398822 -5146
rect 398266 -5702 398502 -5466
rect 398586 -5702 398822 -5466
rect 391986 -6342 392222 -6106
rect 392306 -6342 392542 -6106
rect 391986 -6662 392222 -6426
rect 392306 -6662 392542 -6426
rect 404546 706522 404782 706758
rect 404866 706522 405102 706758
rect 404546 706202 404782 706438
rect 404866 706202 405102 706438
rect 404546 690938 404782 691174
rect 404866 690938 405102 691174
rect 404546 690618 404782 690854
rect 404866 690618 405102 690854
rect 404546 654938 404782 655174
rect 404866 654938 405102 655174
rect 404546 654618 404782 654854
rect 404866 654618 405102 654854
rect 404546 618938 404782 619174
rect 404866 618938 405102 619174
rect 404546 618618 404782 618854
rect 404866 618618 405102 618854
rect 404546 582938 404782 583174
rect 404866 582938 405102 583174
rect 404546 582618 404782 582854
rect 404866 582618 405102 582854
rect 404546 546938 404782 547174
rect 404866 546938 405102 547174
rect 404546 546618 404782 546854
rect 404866 546618 405102 546854
rect 404546 510938 404782 511174
rect 404866 510938 405102 511174
rect 404546 510618 404782 510854
rect 404866 510618 405102 510854
rect 404546 474938 404782 475174
rect 404866 474938 405102 475174
rect 404546 474618 404782 474854
rect 404866 474618 405102 474854
rect 404546 438938 404782 439174
rect 404866 438938 405102 439174
rect 404546 438618 404782 438854
rect 404866 438618 405102 438854
rect 404546 402938 404782 403174
rect 404866 402938 405102 403174
rect 404546 402618 404782 402854
rect 404866 402618 405102 402854
rect 404546 366938 404782 367174
rect 404866 366938 405102 367174
rect 404546 366618 404782 366854
rect 404866 366618 405102 366854
rect 404546 330938 404782 331174
rect 404866 330938 405102 331174
rect 404546 330618 404782 330854
rect 404866 330618 405102 330854
rect 404546 294938 404782 295174
rect 404866 294938 405102 295174
rect 404546 294618 404782 294854
rect 404866 294618 405102 294854
rect 404546 258938 404782 259174
rect 404866 258938 405102 259174
rect 404546 258618 404782 258854
rect 404866 258618 405102 258854
rect 404546 222938 404782 223174
rect 404866 222938 405102 223174
rect 404546 222618 404782 222854
rect 404866 222618 405102 222854
rect 404546 186938 404782 187174
rect 404866 186938 405102 187174
rect 404546 186618 404782 186854
rect 404866 186618 405102 186854
rect 404546 150938 404782 151174
rect 404866 150938 405102 151174
rect 404546 150618 404782 150854
rect 404866 150618 405102 150854
rect 404546 114938 404782 115174
rect 404866 114938 405102 115174
rect 404546 114618 404782 114854
rect 404866 114618 405102 114854
rect 404546 78938 404782 79174
rect 404866 78938 405102 79174
rect 404546 78618 404782 78854
rect 404866 78618 405102 78854
rect 404546 42938 404782 43174
rect 404866 42938 405102 43174
rect 404546 42618 404782 42854
rect 404866 42618 405102 42854
rect 404546 6938 404782 7174
rect 404866 6938 405102 7174
rect 404546 6618 404782 6854
rect 404866 6618 405102 6854
rect 404546 -2502 404782 -2266
rect 404866 -2502 405102 -2266
rect 404546 -2822 404782 -2586
rect 404866 -2822 405102 -2586
rect 408266 694658 408502 694894
rect 408586 694658 408822 694894
rect 408266 694338 408502 694574
rect 408586 694338 408822 694574
rect 408266 658658 408502 658894
rect 408586 658658 408822 658894
rect 408266 658338 408502 658574
rect 408586 658338 408822 658574
rect 408266 622658 408502 622894
rect 408586 622658 408822 622894
rect 408266 622338 408502 622574
rect 408586 622338 408822 622574
rect 408266 586658 408502 586894
rect 408586 586658 408822 586894
rect 408266 586338 408502 586574
rect 408586 586338 408822 586574
rect 408266 550658 408502 550894
rect 408586 550658 408822 550894
rect 408266 550338 408502 550574
rect 408586 550338 408822 550574
rect 408266 514658 408502 514894
rect 408586 514658 408822 514894
rect 408266 514338 408502 514574
rect 408586 514338 408822 514574
rect 408266 478658 408502 478894
rect 408586 478658 408822 478894
rect 408266 478338 408502 478574
rect 408586 478338 408822 478574
rect 408266 442658 408502 442894
rect 408586 442658 408822 442894
rect 408266 442338 408502 442574
rect 408586 442338 408822 442574
rect 408266 406658 408502 406894
rect 408586 406658 408822 406894
rect 408266 406338 408502 406574
rect 408586 406338 408822 406574
rect 408266 370658 408502 370894
rect 408586 370658 408822 370894
rect 408266 370338 408502 370574
rect 408586 370338 408822 370574
rect 408266 334658 408502 334894
rect 408586 334658 408822 334894
rect 408266 334338 408502 334574
rect 408586 334338 408822 334574
rect 408266 298658 408502 298894
rect 408586 298658 408822 298894
rect 408266 298338 408502 298574
rect 408586 298338 408822 298574
rect 408266 262658 408502 262894
rect 408586 262658 408822 262894
rect 408266 262338 408502 262574
rect 408586 262338 408822 262574
rect 408266 226658 408502 226894
rect 408586 226658 408822 226894
rect 408266 226338 408502 226574
rect 408586 226338 408822 226574
rect 408266 190658 408502 190894
rect 408586 190658 408822 190894
rect 408266 190338 408502 190574
rect 408586 190338 408822 190574
rect 408266 154658 408502 154894
rect 408586 154658 408822 154894
rect 408266 154338 408502 154574
rect 408586 154338 408822 154574
rect 408266 118658 408502 118894
rect 408586 118658 408822 118894
rect 408266 118338 408502 118574
rect 408586 118338 408822 118574
rect 408266 82658 408502 82894
rect 408586 82658 408822 82894
rect 408266 82338 408502 82574
rect 408586 82338 408822 82574
rect 408266 46658 408502 46894
rect 408586 46658 408822 46894
rect 408266 46338 408502 46574
rect 408586 46338 408822 46574
rect 408266 10658 408502 10894
rect 408586 10658 408822 10894
rect 408266 10338 408502 10574
rect 408586 10338 408822 10574
rect 410826 705562 411062 705798
rect 411146 705562 411382 705798
rect 410826 705242 411062 705478
rect 411146 705242 411382 705478
rect 410826 669218 411062 669454
rect 411146 669218 411382 669454
rect 410826 668898 411062 669134
rect 411146 668898 411382 669134
rect 410826 633218 411062 633454
rect 411146 633218 411382 633454
rect 410826 632898 411062 633134
rect 411146 632898 411382 633134
rect 410826 597218 411062 597454
rect 411146 597218 411382 597454
rect 410826 596898 411062 597134
rect 411146 596898 411382 597134
rect 410826 561218 411062 561454
rect 411146 561218 411382 561454
rect 410826 560898 411062 561134
rect 411146 560898 411382 561134
rect 410826 525218 411062 525454
rect 411146 525218 411382 525454
rect 410826 524898 411062 525134
rect 411146 524898 411382 525134
rect 410826 489218 411062 489454
rect 411146 489218 411382 489454
rect 410826 488898 411062 489134
rect 411146 488898 411382 489134
rect 410826 453218 411062 453454
rect 411146 453218 411382 453454
rect 410826 452898 411062 453134
rect 411146 452898 411382 453134
rect 410826 417218 411062 417454
rect 411146 417218 411382 417454
rect 410826 416898 411062 417134
rect 411146 416898 411382 417134
rect 410826 381218 411062 381454
rect 411146 381218 411382 381454
rect 410826 380898 411062 381134
rect 411146 380898 411382 381134
rect 410826 345218 411062 345454
rect 411146 345218 411382 345454
rect 410826 344898 411062 345134
rect 411146 344898 411382 345134
rect 410826 309218 411062 309454
rect 411146 309218 411382 309454
rect 410826 308898 411062 309134
rect 411146 308898 411382 309134
rect 410826 273218 411062 273454
rect 411146 273218 411382 273454
rect 410826 272898 411062 273134
rect 411146 272898 411382 273134
rect 410826 237218 411062 237454
rect 411146 237218 411382 237454
rect 410826 236898 411062 237134
rect 411146 236898 411382 237134
rect 410826 201218 411062 201454
rect 411146 201218 411382 201454
rect 410826 200898 411062 201134
rect 411146 200898 411382 201134
rect 410826 165218 411062 165454
rect 411146 165218 411382 165454
rect 410826 164898 411062 165134
rect 411146 164898 411382 165134
rect 410826 129218 411062 129454
rect 411146 129218 411382 129454
rect 410826 128898 411062 129134
rect 411146 128898 411382 129134
rect 410826 93218 411062 93454
rect 411146 93218 411382 93454
rect 410826 92898 411062 93134
rect 411146 92898 411382 93134
rect 410826 57218 411062 57454
rect 411146 57218 411382 57454
rect 410826 56898 411062 57134
rect 411146 56898 411382 57134
rect 410826 21218 411062 21454
rect 411146 21218 411382 21454
rect 410826 20898 411062 21134
rect 411146 20898 411382 21134
rect 410826 -1542 411062 -1306
rect 411146 -1542 411382 -1306
rect 410826 -1862 411062 -1626
rect 411146 -1862 411382 -1626
rect 421986 711322 422222 711558
rect 422306 711322 422542 711558
rect 421986 711002 422222 711238
rect 422306 711002 422542 711238
rect 418266 709402 418502 709638
rect 418586 709402 418822 709638
rect 418266 709082 418502 709318
rect 418586 709082 418822 709318
rect 411986 698378 412222 698614
rect 412306 698378 412542 698614
rect 411986 698058 412222 698294
rect 412306 698058 412542 698294
rect 411986 662378 412222 662614
rect 412306 662378 412542 662614
rect 411986 662058 412222 662294
rect 412306 662058 412542 662294
rect 411986 626378 412222 626614
rect 412306 626378 412542 626614
rect 411986 626058 412222 626294
rect 412306 626058 412542 626294
rect 411986 590378 412222 590614
rect 412306 590378 412542 590614
rect 411986 590058 412222 590294
rect 412306 590058 412542 590294
rect 411986 554378 412222 554614
rect 412306 554378 412542 554614
rect 411986 554058 412222 554294
rect 412306 554058 412542 554294
rect 411986 518378 412222 518614
rect 412306 518378 412542 518614
rect 411986 518058 412222 518294
rect 412306 518058 412542 518294
rect 411986 482378 412222 482614
rect 412306 482378 412542 482614
rect 411986 482058 412222 482294
rect 412306 482058 412542 482294
rect 411986 446378 412222 446614
rect 412306 446378 412542 446614
rect 411986 446058 412222 446294
rect 412306 446058 412542 446294
rect 411986 410378 412222 410614
rect 412306 410378 412542 410614
rect 411986 410058 412222 410294
rect 412306 410058 412542 410294
rect 411986 374378 412222 374614
rect 412306 374378 412542 374614
rect 411986 374058 412222 374294
rect 412306 374058 412542 374294
rect 411986 338378 412222 338614
rect 412306 338378 412542 338614
rect 411986 338058 412222 338294
rect 412306 338058 412542 338294
rect 411986 302378 412222 302614
rect 412306 302378 412542 302614
rect 411986 302058 412222 302294
rect 412306 302058 412542 302294
rect 411986 266378 412222 266614
rect 412306 266378 412542 266614
rect 411986 266058 412222 266294
rect 412306 266058 412542 266294
rect 411986 230378 412222 230614
rect 412306 230378 412542 230614
rect 411986 230058 412222 230294
rect 412306 230058 412542 230294
rect 411986 194378 412222 194614
rect 412306 194378 412542 194614
rect 411986 194058 412222 194294
rect 412306 194058 412542 194294
rect 411986 158378 412222 158614
rect 412306 158378 412542 158614
rect 411986 158058 412222 158294
rect 412306 158058 412542 158294
rect 411986 122378 412222 122614
rect 412306 122378 412542 122614
rect 411986 122058 412222 122294
rect 412306 122058 412542 122294
rect 411986 86378 412222 86614
rect 412306 86378 412542 86614
rect 411986 86058 412222 86294
rect 412306 86058 412542 86294
rect 411986 50378 412222 50614
rect 412306 50378 412542 50614
rect 411986 50058 412222 50294
rect 412306 50058 412542 50294
rect 411986 14378 412222 14614
rect 412306 14378 412542 14614
rect 411986 14058 412222 14294
rect 412306 14058 412542 14294
rect 408266 -4422 408502 -4186
rect 408586 -4422 408822 -4186
rect 408266 -4742 408502 -4506
rect 408586 -4742 408822 -4506
rect 401986 -7302 402222 -7066
rect 402306 -7302 402542 -7066
rect 401986 -7622 402222 -7386
rect 402306 -7622 402542 -7386
rect 414546 707482 414782 707718
rect 414866 707482 415102 707718
rect 414546 707162 414782 707398
rect 414866 707162 415102 707398
rect 414546 672938 414782 673174
rect 414866 672938 415102 673174
rect 414546 672618 414782 672854
rect 414866 672618 415102 672854
rect 414546 636938 414782 637174
rect 414866 636938 415102 637174
rect 414546 636618 414782 636854
rect 414866 636618 415102 636854
rect 414546 600938 414782 601174
rect 414866 600938 415102 601174
rect 414546 600618 414782 600854
rect 414866 600618 415102 600854
rect 414546 564938 414782 565174
rect 414866 564938 415102 565174
rect 414546 564618 414782 564854
rect 414866 564618 415102 564854
rect 414546 528938 414782 529174
rect 414866 528938 415102 529174
rect 414546 528618 414782 528854
rect 414866 528618 415102 528854
rect 414546 492938 414782 493174
rect 414866 492938 415102 493174
rect 414546 492618 414782 492854
rect 414866 492618 415102 492854
rect 414546 456938 414782 457174
rect 414866 456938 415102 457174
rect 414546 456618 414782 456854
rect 414866 456618 415102 456854
rect 414546 420938 414782 421174
rect 414866 420938 415102 421174
rect 414546 420618 414782 420854
rect 414866 420618 415102 420854
rect 414546 384938 414782 385174
rect 414866 384938 415102 385174
rect 414546 384618 414782 384854
rect 414866 384618 415102 384854
rect 414546 348938 414782 349174
rect 414866 348938 415102 349174
rect 414546 348618 414782 348854
rect 414866 348618 415102 348854
rect 414546 312938 414782 313174
rect 414866 312938 415102 313174
rect 414546 312618 414782 312854
rect 414866 312618 415102 312854
rect 414546 276938 414782 277174
rect 414866 276938 415102 277174
rect 414546 276618 414782 276854
rect 414866 276618 415102 276854
rect 414546 240938 414782 241174
rect 414866 240938 415102 241174
rect 414546 240618 414782 240854
rect 414866 240618 415102 240854
rect 414546 204938 414782 205174
rect 414866 204938 415102 205174
rect 414546 204618 414782 204854
rect 414866 204618 415102 204854
rect 414546 168938 414782 169174
rect 414866 168938 415102 169174
rect 414546 168618 414782 168854
rect 414866 168618 415102 168854
rect 414546 132938 414782 133174
rect 414866 132938 415102 133174
rect 414546 132618 414782 132854
rect 414866 132618 415102 132854
rect 414546 96938 414782 97174
rect 414866 96938 415102 97174
rect 414546 96618 414782 96854
rect 414866 96618 415102 96854
rect 414546 60938 414782 61174
rect 414866 60938 415102 61174
rect 414546 60618 414782 60854
rect 414866 60618 415102 60854
rect 414546 24938 414782 25174
rect 414866 24938 415102 25174
rect 414546 24618 414782 24854
rect 414866 24618 415102 24854
rect 414546 -3462 414782 -3226
rect 414866 -3462 415102 -3226
rect 414546 -3782 414782 -3546
rect 414866 -3782 415102 -3546
rect 418266 676658 418502 676894
rect 418586 676658 418822 676894
rect 418266 676338 418502 676574
rect 418586 676338 418822 676574
rect 418266 640658 418502 640894
rect 418586 640658 418822 640894
rect 418266 640338 418502 640574
rect 418586 640338 418822 640574
rect 418266 604658 418502 604894
rect 418586 604658 418822 604894
rect 418266 604338 418502 604574
rect 418586 604338 418822 604574
rect 418266 568658 418502 568894
rect 418586 568658 418822 568894
rect 418266 568338 418502 568574
rect 418586 568338 418822 568574
rect 418266 532658 418502 532894
rect 418586 532658 418822 532894
rect 418266 532338 418502 532574
rect 418586 532338 418822 532574
rect 418266 496658 418502 496894
rect 418586 496658 418822 496894
rect 418266 496338 418502 496574
rect 418586 496338 418822 496574
rect 418266 460658 418502 460894
rect 418586 460658 418822 460894
rect 418266 460338 418502 460574
rect 418586 460338 418822 460574
rect 418266 424658 418502 424894
rect 418586 424658 418822 424894
rect 418266 424338 418502 424574
rect 418586 424338 418822 424574
rect 418266 388658 418502 388894
rect 418586 388658 418822 388894
rect 418266 388338 418502 388574
rect 418586 388338 418822 388574
rect 418266 352658 418502 352894
rect 418586 352658 418822 352894
rect 418266 352338 418502 352574
rect 418586 352338 418822 352574
rect 418266 316658 418502 316894
rect 418586 316658 418822 316894
rect 418266 316338 418502 316574
rect 418586 316338 418822 316574
rect 418266 280658 418502 280894
rect 418586 280658 418822 280894
rect 418266 280338 418502 280574
rect 418586 280338 418822 280574
rect 418266 244658 418502 244894
rect 418586 244658 418822 244894
rect 418266 244338 418502 244574
rect 418586 244338 418822 244574
rect 418266 208658 418502 208894
rect 418586 208658 418822 208894
rect 418266 208338 418502 208574
rect 418586 208338 418822 208574
rect 418266 172658 418502 172894
rect 418586 172658 418822 172894
rect 418266 172338 418502 172574
rect 418586 172338 418822 172574
rect 418266 136658 418502 136894
rect 418586 136658 418822 136894
rect 418266 136338 418502 136574
rect 418586 136338 418822 136574
rect 418266 100658 418502 100894
rect 418586 100658 418822 100894
rect 418266 100338 418502 100574
rect 418586 100338 418822 100574
rect 418266 64658 418502 64894
rect 418586 64658 418822 64894
rect 418266 64338 418502 64574
rect 418586 64338 418822 64574
rect 418266 28658 418502 28894
rect 418586 28658 418822 28894
rect 418266 28338 418502 28574
rect 418586 28338 418822 28574
rect 420826 704602 421062 704838
rect 421146 704602 421382 704838
rect 420826 704282 421062 704518
rect 421146 704282 421382 704518
rect 420826 687218 421062 687454
rect 421146 687218 421382 687454
rect 420826 686898 421062 687134
rect 421146 686898 421382 687134
rect 420826 651218 421062 651454
rect 421146 651218 421382 651454
rect 420826 650898 421062 651134
rect 421146 650898 421382 651134
rect 420826 615218 421062 615454
rect 421146 615218 421382 615454
rect 420826 614898 421062 615134
rect 421146 614898 421382 615134
rect 420826 579218 421062 579454
rect 421146 579218 421382 579454
rect 420826 578898 421062 579134
rect 421146 578898 421382 579134
rect 420826 543218 421062 543454
rect 421146 543218 421382 543454
rect 420826 542898 421062 543134
rect 421146 542898 421382 543134
rect 420826 507218 421062 507454
rect 421146 507218 421382 507454
rect 420826 506898 421062 507134
rect 421146 506898 421382 507134
rect 420826 471218 421062 471454
rect 421146 471218 421382 471454
rect 420826 470898 421062 471134
rect 421146 470898 421382 471134
rect 420826 435218 421062 435454
rect 421146 435218 421382 435454
rect 420826 434898 421062 435134
rect 421146 434898 421382 435134
rect 420826 399218 421062 399454
rect 421146 399218 421382 399454
rect 420826 398898 421062 399134
rect 421146 398898 421382 399134
rect 420826 363218 421062 363454
rect 421146 363218 421382 363454
rect 420826 362898 421062 363134
rect 421146 362898 421382 363134
rect 420826 327218 421062 327454
rect 421146 327218 421382 327454
rect 420826 326898 421062 327134
rect 421146 326898 421382 327134
rect 420826 291218 421062 291454
rect 421146 291218 421382 291454
rect 420826 290898 421062 291134
rect 421146 290898 421382 291134
rect 420826 255218 421062 255454
rect 421146 255218 421382 255454
rect 420826 254898 421062 255134
rect 421146 254898 421382 255134
rect 420826 219218 421062 219454
rect 421146 219218 421382 219454
rect 420826 218898 421062 219134
rect 421146 218898 421382 219134
rect 420826 183218 421062 183454
rect 421146 183218 421382 183454
rect 420826 182898 421062 183134
rect 421146 182898 421382 183134
rect 420826 147218 421062 147454
rect 421146 147218 421382 147454
rect 420826 146898 421062 147134
rect 421146 146898 421382 147134
rect 420826 111218 421062 111454
rect 421146 111218 421382 111454
rect 420826 110898 421062 111134
rect 421146 110898 421382 111134
rect 420826 75218 421062 75454
rect 421146 75218 421382 75454
rect 420826 74898 421062 75134
rect 421146 74898 421382 75134
rect 420826 39218 421062 39454
rect 421146 39218 421382 39454
rect 420826 38898 421062 39134
rect 421146 38898 421382 39134
rect 420826 3218 421062 3454
rect 421146 3218 421382 3454
rect 420826 2898 421062 3134
rect 421146 2898 421382 3134
rect 420826 -582 421062 -346
rect 421146 -582 421382 -346
rect 420826 -902 421062 -666
rect 421146 -902 421382 -666
rect 431986 710362 432222 710598
rect 432306 710362 432542 710598
rect 431986 710042 432222 710278
rect 432306 710042 432542 710278
rect 428266 708442 428502 708678
rect 428586 708442 428822 708678
rect 428266 708122 428502 708358
rect 428586 708122 428822 708358
rect 421986 680378 422222 680614
rect 422306 680378 422542 680614
rect 421986 680058 422222 680294
rect 422306 680058 422542 680294
rect 421986 644378 422222 644614
rect 422306 644378 422542 644614
rect 421986 644058 422222 644294
rect 422306 644058 422542 644294
rect 421986 608378 422222 608614
rect 422306 608378 422542 608614
rect 421986 608058 422222 608294
rect 422306 608058 422542 608294
rect 421986 572378 422222 572614
rect 422306 572378 422542 572614
rect 421986 572058 422222 572294
rect 422306 572058 422542 572294
rect 421986 536378 422222 536614
rect 422306 536378 422542 536614
rect 421986 536058 422222 536294
rect 422306 536058 422542 536294
rect 421986 500378 422222 500614
rect 422306 500378 422542 500614
rect 421986 500058 422222 500294
rect 422306 500058 422542 500294
rect 421986 464378 422222 464614
rect 422306 464378 422542 464614
rect 421986 464058 422222 464294
rect 422306 464058 422542 464294
rect 421986 428378 422222 428614
rect 422306 428378 422542 428614
rect 421986 428058 422222 428294
rect 422306 428058 422542 428294
rect 421986 392378 422222 392614
rect 422306 392378 422542 392614
rect 421986 392058 422222 392294
rect 422306 392058 422542 392294
rect 421986 356378 422222 356614
rect 422306 356378 422542 356614
rect 421986 356058 422222 356294
rect 422306 356058 422542 356294
rect 421986 320378 422222 320614
rect 422306 320378 422542 320614
rect 421986 320058 422222 320294
rect 422306 320058 422542 320294
rect 421986 284378 422222 284614
rect 422306 284378 422542 284614
rect 421986 284058 422222 284294
rect 422306 284058 422542 284294
rect 421986 248378 422222 248614
rect 422306 248378 422542 248614
rect 421986 248058 422222 248294
rect 422306 248058 422542 248294
rect 421986 212378 422222 212614
rect 422306 212378 422542 212614
rect 421986 212058 422222 212294
rect 422306 212058 422542 212294
rect 421986 176378 422222 176614
rect 422306 176378 422542 176614
rect 421986 176058 422222 176294
rect 422306 176058 422542 176294
rect 421986 140378 422222 140614
rect 422306 140378 422542 140614
rect 421986 140058 422222 140294
rect 422306 140058 422542 140294
rect 421986 104378 422222 104614
rect 422306 104378 422542 104614
rect 421986 104058 422222 104294
rect 422306 104058 422542 104294
rect 421986 68378 422222 68614
rect 422306 68378 422542 68614
rect 421986 68058 422222 68294
rect 422306 68058 422542 68294
rect 421986 32378 422222 32614
rect 422306 32378 422542 32614
rect 421986 32058 422222 32294
rect 422306 32058 422542 32294
rect 418266 -5382 418502 -5146
rect 418586 -5382 418822 -5146
rect 418266 -5702 418502 -5466
rect 418586 -5702 418822 -5466
rect 411986 -6342 412222 -6106
rect 412306 -6342 412542 -6106
rect 411986 -6662 412222 -6426
rect 412306 -6662 412542 -6426
rect 424546 706522 424782 706758
rect 424866 706522 425102 706758
rect 424546 706202 424782 706438
rect 424866 706202 425102 706438
rect 424546 690938 424782 691174
rect 424866 690938 425102 691174
rect 424546 690618 424782 690854
rect 424866 690618 425102 690854
rect 424546 654938 424782 655174
rect 424866 654938 425102 655174
rect 424546 654618 424782 654854
rect 424866 654618 425102 654854
rect 424546 618938 424782 619174
rect 424866 618938 425102 619174
rect 424546 618618 424782 618854
rect 424866 618618 425102 618854
rect 424546 582938 424782 583174
rect 424866 582938 425102 583174
rect 424546 582618 424782 582854
rect 424866 582618 425102 582854
rect 424546 546938 424782 547174
rect 424866 546938 425102 547174
rect 424546 546618 424782 546854
rect 424866 546618 425102 546854
rect 424546 510938 424782 511174
rect 424866 510938 425102 511174
rect 424546 510618 424782 510854
rect 424866 510618 425102 510854
rect 424546 474938 424782 475174
rect 424866 474938 425102 475174
rect 424546 474618 424782 474854
rect 424866 474618 425102 474854
rect 424546 438938 424782 439174
rect 424866 438938 425102 439174
rect 424546 438618 424782 438854
rect 424866 438618 425102 438854
rect 424546 402938 424782 403174
rect 424866 402938 425102 403174
rect 424546 402618 424782 402854
rect 424866 402618 425102 402854
rect 424546 366938 424782 367174
rect 424866 366938 425102 367174
rect 424546 366618 424782 366854
rect 424866 366618 425102 366854
rect 424546 330938 424782 331174
rect 424866 330938 425102 331174
rect 424546 330618 424782 330854
rect 424866 330618 425102 330854
rect 424546 294938 424782 295174
rect 424866 294938 425102 295174
rect 424546 294618 424782 294854
rect 424866 294618 425102 294854
rect 424546 258938 424782 259174
rect 424866 258938 425102 259174
rect 424546 258618 424782 258854
rect 424866 258618 425102 258854
rect 424546 222938 424782 223174
rect 424866 222938 425102 223174
rect 424546 222618 424782 222854
rect 424866 222618 425102 222854
rect 424546 186938 424782 187174
rect 424866 186938 425102 187174
rect 424546 186618 424782 186854
rect 424866 186618 425102 186854
rect 424546 150938 424782 151174
rect 424866 150938 425102 151174
rect 424546 150618 424782 150854
rect 424866 150618 425102 150854
rect 424546 114938 424782 115174
rect 424866 114938 425102 115174
rect 424546 114618 424782 114854
rect 424866 114618 425102 114854
rect 424546 78938 424782 79174
rect 424866 78938 425102 79174
rect 424546 78618 424782 78854
rect 424866 78618 425102 78854
rect 424546 42938 424782 43174
rect 424866 42938 425102 43174
rect 424546 42618 424782 42854
rect 424866 42618 425102 42854
rect 424546 6938 424782 7174
rect 424866 6938 425102 7174
rect 424546 6618 424782 6854
rect 424866 6618 425102 6854
rect 424546 -2502 424782 -2266
rect 424866 -2502 425102 -2266
rect 424546 -2822 424782 -2586
rect 424866 -2822 425102 -2586
rect 428266 694658 428502 694894
rect 428586 694658 428822 694894
rect 428266 694338 428502 694574
rect 428586 694338 428822 694574
rect 428266 658658 428502 658894
rect 428586 658658 428822 658894
rect 428266 658338 428502 658574
rect 428586 658338 428822 658574
rect 428266 622658 428502 622894
rect 428586 622658 428822 622894
rect 428266 622338 428502 622574
rect 428586 622338 428822 622574
rect 428266 586658 428502 586894
rect 428586 586658 428822 586894
rect 428266 586338 428502 586574
rect 428586 586338 428822 586574
rect 428266 550658 428502 550894
rect 428586 550658 428822 550894
rect 428266 550338 428502 550574
rect 428586 550338 428822 550574
rect 428266 514658 428502 514894
rect 428586 514658 428822 514894
rect 428266 514338 428502 514574
rect 428586 514338 428822 514574
rect 428266 478658 428502 478894
rect 428586 478658 428822 478894
rect 428266 478338 428502 478574
rect 428586 478338 428822 478574
rect 428266 442658 428502 442894
rect 428586 442658 428822 442894
rect 428266 442338 428502 442574
rect 428586 442338 428822 442574
rect 428266 406658 428502 406894
rect 428586 406658 428822 406894
rect 428266 406338 428502 406574
rect 428586 406338 428822 406574
rect 428266 370658 428502 370894
rect 428586 370658 428822 370894
rect 428266 370338 428502 370574
rect 428586 370338 428822 370574
rect 428266 334658 428502 334894
rect 428586 334658 428822 334894
rect 428266 334338 428502 334574
rect 428586 334338 428822 334574
rect 428266 298658 428502 298894
rect 428586 298658 428822 298894
rect 428266 298338 428502 298574
rect 428586 298338 428822 298574
rect 428266 262658 428502 262894
rect 428586 262658 428822 262894
rect 428266 262338 428502 262574
rect 428586 262338 428822 262574
rect 428266 226658 428502 226894
rect 428586 226658 428822 226894
rect 428266 226338 428502 226574
rect 428586 226338 428822 226574
rect 428266 190658 428502 190894
rect 428586 190658 428822 190894
rect 428266 190338 428502 190574
rect 428586 190338 428822 190574
rect 428266 154658 428502 154894
rect 428586 154658 428822 154894
rect 428266 154338 428502 154574
rect 428586 154338 428822 154574
rect 428266 118658 428502 118894
rect 428586 118658 428822 118894
rect 428266 118338 428502 118574
rect 428586 118338 428822 118574
rect 428266 82658 428502 82894
rect 428586 82658 428822 82894
rect 428266 82338 428502 82574
rect 428586 82338 428822 82574
rect 428266 46658 428502 46894
rect 428586 46658 428822 46894
rect 428266 46338 428502 46574
rect 428586 46338 428822 46574
rect 428266 10658 428502 10894
rect 428586 10658 428822 10894
rect 428266 10338 428502 10574
rect 428586 10338 428822 10574
rect 430826 705562 431062 705798
rect 431146 705562 431382 705798
rect 430826 705242 431062 705478
rect 431146 705242 431382 705478
rect 430826 669218 431062 669454
rect 431146 669218 431382 669454
rect 430826 668898 431062 669134
rect 431146 668898 431382 669134
rect 430826 633218 431062 633454
rect 431146 633218 431382 633454
rect 430826 632898 431062 633134
rect 431146 632898 431382 633134
rect 430826 597218 431062 597454
rect 431146 597218 431382 597454
rect 430826 596898 431062 597134
rect 431146 596898 431382 597134
rect 430826 561218 431062 561454
rect 431146 561218 431382 561454
rect 430826 560898 431062 561134
rect 431146 560898 431382 561134
rect 430826 525218 431062 525454
rect 431146 525218 431382 525454
rect 430826 524898 431062 525134
rect 431146 524898 431382 525134
rect 430826 489218 431062 489454
rect 431146 489218 431382 489454
rect 430826 488898 431062 489134
rect 431146 488898 431382 489134
rect 430826 453218 431062 453454
rect 431146 453218 431382 453454
rect 430826 452898 431062 453134
rect 431146 452898 431382 453134
rect 430826 417218 431062 417454
rect 431146 417218 431382 417454
rect 430826 416898 431062 417134
rect 431146 416898 431382 417134
rect 430826 381218 431062 381454
rect 431146 381218 431382 381454
rect 430826 380898 431062 381134
rect 431146 380898 431382 381134
rect 430826 345218 431062 345454
rect 431146 345218 431382 345454
rect 430826 344898 431062 345134
rect 431146 344898 431382 345134
rect 430826 309218 431062 309454
rect 431146 309218 431382 309454
rect 430826 308898 431062 309134
rect 431146 308898 431382 309134
rect 430826 273218 431062 273454
rect 431146 273218 431382 273454
rect 430826 272898 431062 273134
rect 431146 272898 431382 273134
rect 430826 237218 431062 237454
rect 431146 237218 431382 237454
rect 430826 236898 431062 237134
rect 431146 236898 431382 237134
rect 430826 201218 431062 201454
rect 431146 201218 431382 201454
rect 430826 200898 431062 201134
rect 431146 200898 431382 201134
rect 430826 165218 431062 165454
rect 431146 165218 431382 165454
rect 430826 164898 431062 165134
rect 431146 164898 431382 165134
rect 430826 129218 431062 129454
rect 431146 129218 431382 129454
rect 430826 128898 431062 129134
rect 431146 128898 431382 129134
rect 430826 93218 431062 93454
rect 431146 93218 431382 93454
rect 430826 92898 431062 93134
rect 431146 92898 431382 93134
rect 430826 57218 431062 57454
rect 431146 57218 431382 57454
rect 430826 56898 431062 57134
rect 431146 56898 431382 57134
rect 430826 21218 431062 21454
rect 431146 21218 431382 21454
rect 430826 20898 431062 21134
rect 431146 20898 431382 21134
rect 430826 -1542 431062 -1306
rect 431146 -1542 431382 -1306
rect 430826 -1862 431062 -1626
rect 431146 -1862 431382 -1626
rect 441986 711322 442222 711558
rect 442306 711322 442542 711558
rect 441986 711002 442222 711238
rect 442306 711002 442542 711238
rect 438266 709402 438502 709638
rect 438586 709402 438822 709638
rect 438266 709082 438502 709318
rect 438586 709082 438822 709318
rect 431986 698378 432222 698614
rect 432306 698378 432542 698614
rect 431986 698058 432222 698294
rect 432306 698058 432542 698294
rect 431986 662378 432222 662614
rect 432306 662378 432542 662614
rect 431986 662058 432222 662294
rect 432306 662058 432542 662294
rect 431986 626378 432222 626614
rect 432306 626378 432542 626614
rect 431986 626058 432222 626294
rect 432306 626058 432542 626294
rect 431986 590378 432222 590614
rect 432306 590378 432542 590614
rect 431986 590058 432222 590294
rect 432306 590058 432542 590294
rect 431986 554378 432222 554614
rect 432306 554378 432542 554614
rect 431986 554058 432222 554294
rect 432306 554058 432542 554294
rect 431986 518378 432222 518614
rect 432306 518378 432542 518614
rect 431986 518058 432222 518294
rect 432306 518058 432542 518294
rect 431986 482378 432222 482614
rect 432306 482378 432542 482614
rect 431986 482058 432222 482294
rect 432306 482058 432542 482294
rect 431986 446378 432222 446614
rect 432306 446378 432542 446614
rect 431986 446058 432222 446294
rect 432306 446058 432542 446294
rect 431986 410378 432222 410614
rect 432306 410378 432542 410614
rect 431986 410058 432222 410294
rect 432306 410058 432542 410294
rect 431986 374378 432222 374614
rect 432306 374378 432542 374614
rect 431986 374058 432222 374294
rect 432306 374058 432542 374294
rect 431986 338378 432222 338614
rect 432306 338378 432542 338614
rect 431986 338058 432222 338294
rect 432306 338058 432542 338294
rect 431986 302378 432222 302614
rect 432306 302378 432542 302614
rect 431986 302058 432222 302294
rect 432306 302058 432542 302294
rect 431986 266378 432222 266614
rect 432306 266378 432542 266614
rect 431986 266058 432222 266294
rect 432306 266058 432542 266294
rect 431986 230378 432222 230614
rect 432306 230378 432542 230614
rect 431986 230058 432222 230294
rect 432306 230058 432542 230294
rect 431986 194378 432222 194614
rect 432306 194378 432542 194614
rect 431986 194058 432222 194294
rect 432306 194058 432542 194294
rect 431986 158378 432222 158614
rect 432306 158378 432542 158614
rect 431986 158058 432222 158294
rect 432306 158058 432542 158294
rect 431986 122378 432222 122614
rect 432306 122378 432542 122614
rect 431986 122058 432222 122294
rect 432306 122058 432542 122294
rect 431986 86378 432222 86614
rect 432306 86378 432542 86614
rect 431986 86058 432222 86294
rect 432306 86058 432542 86294
rect 431986 50378 432222 50614
rect 432306 50378 432542 50614
rect 431986 50058 432222 50294
rect 432306 50058 432542 50294
rect 431986 14378 432222 14614
rect 432306 14378 432542 14614
rect 431986 14058 432222 14294
rect 432306 14058 432542 14294
rect 428266 -4422 428502 -4186
rect 428586 -4422 428822 -4186
rect 428266 -4742 428502 -4506
rect 428586 -4742 428822 -4506
rect 421986 -7302 422222 -7066
rect 422306 -7302 422542 -7066
rect 421986 -7622 422222 -7386
rect 422306 -7622 422542 -7386
rect 434546 707482 434782 707718
rect 434866 707482 435102 707718
rect 434546 707162 434782 707398
rect 434866 707162 435102 707398
rect 434546 672938 434782 673174
rect 434866 672938 435102 673174
rect 434546 672618 434782 672854
rect 434866 672618 435102 672854
rect 434546 636938 434782 637174
rect 434866 636938 435102 637174
rect 434546 636618 434782 636854
rect 434866 636618 435102 636854
rect 434546 600938 434782 601174
rect 434866 600938 435102 601174
rect 434546 600618 434782 600854
rect 434866 600618 435102 600854
rect 434546 564938 434782 565174
rect 434866 564938 435102 565174
rect 434546 564618 434782 564854
rect 434866 564618 435102 564854
rect 434546 528938 434782 529174
rect 434866 528938 435102 529174
rect 434546 528618 434782 528854
rect 434866 528618 435102 528854
rect 434546 492938 434782 493174
rect 434866 492938 435102 493174
rect 434546 492618 434782 492854
rect 434866 492618 435102 492854
rect 434546 456938 434782 457174
rect 434866 456938 435102 457174
rect 434546 456618 434782 456854
rect 434866 456618 435102 456854
rect 434546 420938 434782 421174
rect 434866 420938 435102 421174
rect 434546 420618 434782 420854
rect 434866 420618 435102 420854
rect 434546 384938 434782 385174
rect 434866 384938 435102 385174
rect 434546 384618 434782 384854
rect 434866 384618 435102 384854
rect 434546 348938 434782 349174
rect 434866 348938 435102 349174
rect 434546 348618 434782 348854
rect 434866 348618 435102 348854
rect 434546 312938 434782 313174
rect 434866 312938 435102 313174
rect 434546 312618 434782 312854
rect 434866 312618 435102 312854
rect 434546 276938 434782 277174
rect 434866 276938 435102 277174
rect 434546 276618 434782 276854
rect 434866 276618 435102 276854
rect 434546 240938 434782 241174
rect 434866 240938 435102 241174
rect 434546 240618 434782 240854
rect 434866 240618 435102 240854
rect 434546 204938 434782 205174
rect 434866 204938 435102 205174
rect 434546 204618 434782 204854
rect 434866 204618 435102 204854
rect 434546 168938 434782 169174
rect 434866 168938 435102 169174
rect 434546 168618 434782 168854
rect 434866 168618 435102 168854
rect 434546 132938 434782 133174
rect 434866 132938 435102 133174
rect 434546 132618 434782 132854
rect 434866 132618 435102 132854
rect 434546 96938 434782 97174
rect 434866 96938 435102 97174
rect 434546 96618 434782 96854
rect 434866 96618 435102 96854
rect 434546 60938 434782 61174
rect 434866 60938 435102 61174
rect 434546 60618 434782 60854
rect 434866 60618 435102 60854
rect 434546 24938 434782 25174
rect 434866 24938 435102 25174
rect 434546 24618 434782 24854
rect 434866 24618 435102 24854
rect 434546 -3462 434782 -3226
rect 434866 -3462 435102 -3226
rect 434546 -3782 434782 -3546
rect 434866 -3782 435102 -3546
rect 438266 676658 438502 676894
rect 438586 676658 438822 676894
rect 438266 676338 438502 676574
rect 438586 676338 438822 676574
rect 438266 640658 438502 640894
rect 438586 640658 438822 640894
rect 438266 640338 438502 640574
rect 438586 640338 438822 640574
rect 438266 604658 438502 604894
rect 438586 604658 438822 604894
rect 438266 604338 438502 604574
rect 438586 604338 438822 604574
rect 438266 568658 438502 568894
rect 438586 568658 438822 568894
rect 438266 568338 438502 568574
rect 438586 568338 438822 568574
rect 438266 532658 438502 532894
rect 438586 532658 438822 532894
rect 438266 532338 438502 532574
rect 438586 532338 438822 532574
rect 438266 496658 438502 496894
rect 438586 496658 438822 496894
rect 438266 496338 438502 496574
rect 438586 496338 438822 496574
rect 438266 460658 438502 460894
rect 438586 460658 438822 460894
rect 438266 460338 438502 460574
rect 438586 460338 438822 460574
rect 438266 424658 438502 424894
rect 438586 424658 438822 424894
rect 438266 424338 438502 424574
rect 438586 424338 438822 424574
rect 438266 388658 438502 388894
rect 438586 388658 438822 388894
rect 438266 388338 438502 388574
rect 438586 388338 438822 388574
rect 438266 352658 438502 352894
rect 438586 352658 438822 352894
rect 438266 352338 438502 352574
rect 438586 352338 438822 352574
rect 438266 316658 438502 316894
rect 438586 316658 438822 316894
rect 438266 316338 438502 316574
rect 438586 316338 438822 316574
rect 438266 280658 438502 280894
rect 438586 280658 438822 280894
rect 438266 280338 438502 280574
rect 438586 280338 438822 280574
rect 438266 244658 438502 244894
rect 438586 244658 438822 244894
rect 438266 244338 438502 244574
rect 438586 244338 438822 244574
rect 438266 208658 438502 208894
rect 438586 208658 438822 208894
rect 438266 208338 438502 208574
rect 438586 208338 438822 208574
rect 438266 172658 438502 172894
rect 438586 172658 438822 172894
rect 438266 172338 438502 172574
rect 438586 172338 438822 172574
rect 438266 136658 438502 136894
rect 438586 136658 438822 136894
rect 438266 136338 438502 136574
rect 438586 136338 438822 136574
rect 438266 100658 438502 100894
rect 438586 100658 438822 100894
rect 438266 100338 438502 100574
rect 438586 100338 438822 100574
rect 438266 64658 438502 64894
rect 438586 64658 438822 64894
rect 438266 64338 438502 64574
rect 438586 64338 438822 64574
rect 438266 28658 438502 28894
rect 438586 28658 438822 28894
rect 438266 28338 438502 28574
rect 438586 28338 438822 28574
rect 440826 704602 441062 704838
rect 441146 704602 441382 704838
rect 440826 704282 441062 704518
rect 441146 704282 441382 704518
rect 440826 687218 441062 687454
rect 441146 687218 441382 687454
rect 440826 686898 441062 687134
rect 441146 686898 441382 687134
rect 440826 651218 441062 651454
rect 441146 651218 441382 651454
rect 440826 650898 441062 651134
rect 441146 650898 441382 651134
rect 440826 615218 441062 615454
rect 441146 615218 441382 615454
rect 440826 614898 441062 615134
rect 441146 614898 441382 615134
rect 440826 579218 441062 579454
rect 441146 579218 441382 579454
rect 440826 578898 441062 579134
rect 441146 578898 441382 579134
rect 440826 543218 441062 543454
rect 441146 543218 441382 543454
rect 440826 542898 441062 543134
rect 441146 542898 441382 543134
rect 440826 507218 441062 507454
rect 441146 507218 441382 507454
rect 440826 506898 441062 507134
rect 441146 506898 441382 507134
rect 440826 471218 441062 471454
rect 441146 471218 441382 471454
rect 440826 470898 441062 471134
rect 441146 470898 441382 471134
rect 440826 435218 441062 435454
rect 441146 435218 441382 435454
rect 440826 434898 441062 435134
rect 441146 434898 441382 435134
rect 440826 399218 441062 399454
rect 441146 399218 441382 399454
rect 440826 398898 441062 399134
rect 441146 398898 441382 399134
rect 440826 363218 441062 363454
rect 441146 363218 441382 363454
rect 440826 362898 441062 363134
rect 441146 362898 441382 363134
rect 440826 327218 441062 327454
rect 441146 327218 441382 327454
rect 440826 326898 441062 327134
rect 441146 326898 441382 327134
rect 440826 291218 441062 291454
rect 441146 291218 441382 291454
rect 440826 290898 441062 291134
rect 441146 290898 441382 291134
rect 440826 255218 441062 255454
rect 441146 255218 441382 255454
rect 440826 254898 441062 255134
rect 441146 254898 441382 255134
rect 440826 219218 441062 219454
rect 441146 219218 441382 219454
rect 440826 218898 441062 219134
rect 441146 218898 441382 219134
rect 440826 183218 441062 183454
rect 441146 183218 441382 183454
rect 440826 182898 441062 183134
rect 441146 182898 441382 183134
rect 440826 147218 441062 147454
rect 441146 147218 441382 147454
rect 440826 146898 441062 147134
rect 441146 146898 441382 147134
rect 440826 111218 441062 111454
rect 441146 111218 441382 111454
rect 440826 110898 441062 111134
rect 441146 110898 441382 111134
rect 440826 75218 441062 75454
rect 441146 75218 441382 75454
rect 440826 74898 441062 75134
rect 441146 74898 441382 75134
rect 440826 39218 441062 39454
rect 441146 39218 441382 39454
rect 440826 38898 441062 39134
rect 441146 38898 441382 39134
rect 440826 3218 441062 3454
rect 441146 3218 441382 3454
rect 440826 2898 441062 3134
rect 441146 2898 441382 3134
rect 440826 -582 441062 -346
rect 441146 -582 441382 -346
rect 440826 -902 441062 -666
rect 441146 -902 441382 -666
rect 451986 710362 452222 710598
rect 452306 710362 452542 710598
rect 451986 710042 452222 710278
rect 452306 710042 452542 710278
rect 448266 708442 448502 708678
rect 448586 708442 448822 708678
rect 448266 708122 448502 708358
rect 448586 708122 448822 708358
rect 441986 680378 442222 680614
rect 442306 680378 442542 680614
rect 441986 680058 442222 680294
rect 442306 680058 442542 680294
rect 441986 644378 442222 644614
rect 442306 644378 442542 644614
rect 441986 644058 442222 644294
rect 442306 644058 442542 644294
rect 441986 608378 442222 608614
rect 442306 608378 442542 608614
rect 441986 608058 442222 608294
rect 442306 608058 442542 608294
rect 441986 572378 442222 572614
rect 442306 572378 442542 572614
rect 441986 572058 442222 572294
rect 442306 572058 442542 572294
rect 441986 536378 442222 536614
rect 442306 536378 442542 536614
rect 441986 536058 442222 536294
rect 442306 536058 442542 536294
rect 441986 500378 442222 500614
rect 442306 500378 442542 500614
rect 441986 500058 442222 500294
rect 442306 500058 442542 500294
rect 441986 464378 442222 464614
rect 442306 464378 442542 464614
rect 441986 464058 442222 464294
rect 442306 464058 442542 464294
rect 441986 428378 442222 428614
rect 442306 428378 442542 428614
rect 441986 428058 442222 428294
rect 442306 428058 442542 428294
rect 441986 392378 442222 392614
rect 442306 392378 442542 392614
rect 441986 392058 442222 392294
rect 442306 392058 442542 392294
rect 441986 356378 442222 356614
rect 442306 356378 442542 356614
rect 441986 356058 442222 356294
rect 442306 356058 442542 356294
rect 441986 320378 442222 320614
rect 442306 320378 442542 320614
rect 441986 320058 442222 320294
rect 442306 320058 442542 320294
rect 441986 284378 442222 284614
rect 442306 284378 442542 284614
rect 441986 284058 442222 284294
rect 442306 284058 442542 284294
rect 441986 248378 442222 248614
rect 442306 248378 442542 248614
rect 441986 248058 442222 248294
rect 442306 248058 442542 248294
rect 441986 212378 442222 212614
rect 442306 212378 442542 212614
rect 441986 212058 442222 212294
rect 442306 212058 442542 212294
rect 441986 176378 442222 176614
rect 442306 176378 442542 176614
rect 441986 176058 442222 176294
rect 442306 176058 442542 176294
rect 441986 140378 442222 140614
rect 442306 140378 442542 140614
rect 441986 140058 442222 140294
rect 442306 140058 442542 140294
rect 441986 104378 442222 104614
rect 442306 104378 442542 104614
rect 441986 104058 442222 104294
rect 442306 104058 442542 104294
rect 441986 68378 442222 68614
rect 442306 68378 442542 68614
rect 441986 68058 442222 68294
rect 442306 68058 442542 68294
rect 441986 32378 442222 32614
rect 442306 32378 442542 32614
rect 441986 32058 442222 32294
rect 442306 32058 442542 32294
rect 438266 -5382 438502 -5146
rect 438586 -5382 438822 -5146
rect 438266 -5702 438502 -5466
rect 438586 -5702 438822 -5466
rect 431986 -6342 432222 -6106
rect 432306 -6342 432542 -6106
rect 431986 -6662 432222 -6426
rect 432306 -6662 432542 -6426
rect 444546 706522 444782 706758
rect 444866 706522 445102 706758
rect 444546 706202 444782 706438
rect 444866 706202 445102 706438
rect 444546 690938 444782 691174
rect 444866 690938 445102 691174
rect 444546 690618 444782 690854
rect 444866 690618 445102 690854
rect 444546 654938 444782 655174
rect 444866 654938 445102 655174
rect 444546 654618 444782 654854
rect 444866 654618 445102 654854
rect 444546 618938 444782 619174
rect 444866 618938 445102 619174
rect 444546 618618 444782 618854
rect 444866 618618 445102 618854
rect 444546 582938 444782 583174
rect 444866 582938 445102 583174
rect 444546 582618 444782 582854
rect 444866 582618 445102 582854
rect 444546 546938 444782 547174
rect 444866 546938 445102 547174
rect 444546 546618 444782 546854
rect 444866 546618 445102 546854
rect 444546 510938 444782 511174
rect 444866 510938 445102 511174
rect 444546 510618 444782 510854
rect 444866 510618 445102 510854
rect 444546 474938 444782 475174
rect 444866 474938 445102 475174
rect 444546 474618 444782 474854
rect 444866 474618 445102 474854
rect 444546 438938 444782 439174
rect 444866 438938 445102 439174
rect 444546 438618 444782 438854
rect 444866 438618 445102 438854
rect 444546 402938 444782 403174
rect 444866 402938 445102 403174
rect 444546 402618 444782 402854
rect 444866 402618 445102 402854
rect 444546 366938 444782 367174
rect 444866 366938 445102 367174
rect 444546 366618 444782 366854
rect 444866 366618 445102 366854
rect 444546 330938 444782 331174
rect 444866 330938 445102 331174
rect 444546 330618 444782 330854
rect 444866 330618 445102 330854
rect 444546 294938 444782 295174
rect 444866 294938 445102 295174
rect 444546 294618 444782 294854
rect 444866 294618 445102 294854
rect 444546 258938 444782 259174
rect 444866 258938 445102 259174
rect 444546 258618 444782 258854
rect 444866 258618 445102 258854
rect 444546 222938 444782 223174
rect 444866 222938 445102 223174
rect 444546 222618 444782 222854
rect 444866 222618 445102 222854
rect 444546 186938 444782 187174
rect 444866 186938 445102 187174
rect 444546 186618 444782 186854
rect 444866 186618 445102 186854
rect 444546 150938 444782 151174
rect 444866 150938 445102 151174
rect 444546 150618 444782 150854
rect 444866 150618 445102 150854
rect 444546 114938 444782 115174
rect 444866 114938 445102 115174
rect 444546 114618 444782 114854
rect 444866 114618 445102 114854
rect 444546 78938 444782 79174
rect 444866 78938 445102 79174
rect 444546 78618 444782 78854
rect 444866 78618 445102 78854
rect 444546 42938 444782 43174
rect 444866 42938 445102 43174
rect 444546 42618 444782 42854
rect 444866 42618 445102 42854
rect 444546 6938 444782 7174
rect 444866 6938 445102 7174
rect 444546 6618 444782 6854
rect 444866 6618 445102 6854
rect 444546 -2502 444782 -2266
rect 444866 -2502 445102 -2266
rect 444546 -2822 444782 -2586
rect 444866 -2822 445102 -2586
rect 448266 694658 448502 694894
rect 448586 694658 448822 694894
rect 448266 694338 448502 694574
rect 448586 694338 448822 694574
rect 448266 658658 448502 658894
rect 448586 658658 448822 658894
rect 448266 658338 448502 658574
rect 448586 658338 448822 658574
rect 448266 622658 448502 622894
rect 448586 622658 448822 622894
rect 448266 622338 448502 622574
rect 448586 622338 448822 622574
rect 448266 586658 448502 586894
rect 448586 586658 448822 586894
rect 448266 586338 448502 586574
rect 448586 586338 448822 586574
rect 448266 550658 448502 550894
rect 448586 550658 448822 550894
rect 448266 550338 448502 550574
rect 448586 550338 448822 550574
rect 448266 514658 448502 514894
rect 448586 514658 448822 514894
rect 448266 514338 448502 514574
rect 448586 514338 448822 514574
rect 448266 478658 448502 478894
rect 448586 478658 448822 478894
rect 448266 478338 448502 478574
rect 448586 478338 448822 478574
rect 448266 442658 448502 442894
rect 448586 442658 448822 442894
rect 448266 442338 448502 442574
rect 448586 442338 448822 442574
rect 448266 406658 448502 406894
rect 448586 406658 448822 406894
rect 448266 406338 448502 406574
rect 448586 406338 448822 406574
rect 448266 370658 448502 370894
rect 448586 370658 448822 370894
rect 448266 370338 448502 370574
rect 448586 370338 448822 370574
rect 448266 334658 448502 334894
rect 448586 334658 448822 334894
rect 448266 334338 448502 334574
rect 448586 334338 448822 334574
rect 448266 298658 448502 298894
rect 448586 298658 448822 298894
rect 448266 298338 448502 298574
rect 448586 298338 448822 298574
rect 448266 262658 448502 262894
rect 448586 262658 448822 262894
rect 448266 262338 448502 262574
rect 448586 262338 448822 262574
rect 448266 226658 448502 226894
rect 448586 226658 448822 226894
rect 448266 226338 448502 226574
rect 448586 226338 448822 226574
rect 448266 190658 448502 190894
rect 448586 190658 448822 190894
rect 448266 190338 448502 190574
rect 448586 190338 448822 190574
rect 448266 154658 448502 154894
rect 448586 154658 448822 154894
rect 448266 154338 448502 154574
rect 448586 154338 448822 154574
rect 448266 118658 448502 118894
rect 448586 118658 448822 118894
rect 448266 118338 448502 118574
rect 448586 118338 448822 118574
rect 448266 82658 448502 82894
rect 448586 82658 448822 82894
rect 448266 82338 448502 82574
rect 448586 82338 448822 82574
rect 448266 46658 448502 46894
rect 448586 46658 448822 46894
rect 448266 46338 448502 46574
rect 448586 46338 448822 46574
rect 448266 10658 448502 10894
rect 448586 10658 448822 10894
rect 448266 10338 448502 10574
rect 448586 10338 448822 10574
rect 450826 705562 451062 705798
rect 451146 705562 451382 705798
rect 450826 705242 451062 705478
rect 451146 705242 451382 705478
rect 450826 669218 451062 669454
rect 451146 669218 451382 669454
rect 450826 668898 451062 669134
rect 451146 668898 451382 669134
rect 450826 633218 451062 633454
rect 451146 633218 451382 633454
rect 450826 632898 451062 633134
rect 451146 632898 451382 633134
rect 450826 597218 451062 597454
rect 451146 597218 451382 597454
rect 450826 596898 451062 597134
rect 451146 596898 451382 597134
rect 450826 561218 451062 561454
rect 451146 561218 451382 561454
rect 450826 560898 451062 561134
rect 451146 560898 451382 561134
rect 450826 525218 451062 525454
rect 451146 525218 451382 525454
rect 450826 524898 451062 525134
rect 451146 524898 451382 525134
rect 450826 489218 451062 489454
rect 451146 489218 451382 489454
rect 450826 488898 451062 489134
rect 451146 488898 451382 489134
rect 450826 453218 451062 453454
rect 451146 453218 451382 453454
rect 450826 452898 451062 453134
rect 451146 452898 451382 453134
rect 450826 417218 451062 417454
rect 451146 417218 451382 417454
rect 450826 416898 451062 417134
rect 451146 416898 451382 417134
rect 450826 381218 451062 381454
rect 451146 381218 451382 381454
rect 450826 380898 451062 381134
rect 451146 380898 451382 381134
rect 450826 345218 451062 345454
rect 451146 345218 451382 345454
rect 450826 344898 451062 345134
rect 451146 344898 451382 345134
rect 450826 309218 451062 309454
rect 451146 309218 451382 309454
rect 450826 308898 451062 309134
rect 451146 308898 451382 309134
rect 450826 273218 451062 273454
rect 451146 273218 451382 273454
rect 450826 272898 451062 273134
rect 451146 272898 451382 273134
rect 450826 237218 451062 237454
rect 451146 237218 451382 237454
rect 450826 236898 451062 237134
rect 451146 236898 451382 237134
rect 450826 201218 451062 201454
rect 451146 201218 451382 201454
rect 450826 200898 451062 201134
rect 451146 200898 451382 201134
rect 450826 165218 451062 165454
rect 451146 165218 451382 165454
rect 450826 164898 451062 165134
rect 451146 164898 451382 165134
rect 450826 129218 451062 129454
rect 451146 129218 451382 129454
rect 450826 128898 451062 129134
rect 451146 128898 451382 129134
rect 450826 93218 451062 93454
rect 451146 93218 451382 93454
rect 450826 92898 451062 93134
rect 451146 92898 451382 93134
rect 450826 57218 451062 57454
rect 451146 57218 451382 57454
rect 450826 56898 451062 57134
rect 451146 56898 451382 57134
rect 450826 21218 451062 21454
rect 451146 21218 451382 21454
rect 450826 20898 451062 21134
rect 451146 20898 451382 21134
rect 450826 -1542 451062 -1306
rect 451146 -1542 451382 -1306
rect 450826 -1862 451062 -1626
rect 451146 -1862 451382 -1626
rect 461986 711322 462222 711558
rect 462306 711322 462542 711558
rect 461986 711002 462222 711238
rect 462306 711002 462542 711238
rect 458266 709402 458502 709638
rect 458586 709402 458822 709638
rect 458266 709082 458502 709318
rect 458586 709082 458822 709318
rect 451986 698378 452222 698614
rect 452306 698378 452542 698614
rect 451986 698058 452222 698294
rect 452306 698058 452542 698294
rect 451986 662378 452222 662614
rect 452306 662378 452542 662614
rect 451986 662058 452222 662294
rect 452306 662058 452542 662294
rect 451986 626378 452222 626614
rect 452306 626378 452542 626614
rect 451986 626058 452222 626294
rect 452306 626058 452542 626294
rect 451986 590378 452222 590614
rect 452306 590378 452542 590614
rect 451986 590058 452222 590294
rect 452306 590058 452542 590294
rect 451986 554378 452222 554614
rect 452306 554378 452542 554614
rect 451986 554058 452222 554294
rect 452306 554058 452542 554294
rect 451986 518378 452222 518614
rect 452306 518378 452542 518614
rect 451986 518058 452222 518294
rect 452306 518058 452542 518294
rect 451986 482378 452222 482614
rect 452306 482378 452542 482614
rect 451986 482058 452222 482294
rect 452306 482058 452542 482294
rect 451986 446378 452222 446614
rect 452306 446378 452542 446614
rect 451986 446058 452222 446294
rect 452306 446058 452542 446294
rect 451986 410378 452222 410614
rect 452306 410378 452542 410614
rect 451986 410058 452222 410294
rect 452306 410058 452542 410294
rect 451986 374378 452222 374614
rect 452306 374378 452542 374614
rect 451986 374058 452222 374294
rect 452306 374058 452542 374294
rect 451986 338378 452222 338614
rect 452306 338378 452542 338614
rect 451986 338058 452222 338294
rect 452306 338058 452542 338294
rect 451986 302378 452222 302614
rect 452306 302378 452542 302614
rect 451986 302058 452222 302294
rect 452306 302058 452542 302294
rect 451986 266378 452222 266614
rect 452306 266378 452542 266614
rect 451986 266058 452222 266294
rect 452306 266058 452542 266294
rect 451986 230378 452222 230614
rect 452306 230378 452542 230614
rect 451986 230058 452222 230294
rect 452306 230058 452542 230294
rect 451986 194378 452222 194614
rect 452306 194378 452542 194614
rect 451986 194058 452222 194294
rect 452306 194058 452542 194294
rect 451986 158378 452222 158614
rect 452306 158378 452542 158614
rect 451986 158058 452222 158294
rect 452306 158058 452542 158294
rect 451986 122378 452222 122614
rect 452306 122378 452542 122614
rect 451986 122058 452222 122294
rect 452306 122058 452542 122294
rect 451986 86378 452222 86614
rect 452306 86378 452542 86614
rect 451986 86058 452222 86294
rect 452306 86058 452542 86294
rect 451986 50378 452222 50614
rect 452306 50378 452542 50614
rect 451986 50058 452222 50294
rect 452306 50058 452542 50294
rect 451986 14378 452222 14614
rect 452306 14378 452542 14614
rect 451986 14058 452222 14294
rect 452306 14058 452542 14294
rect 448266 -4422 448502 -4186
rect 448586 -4422 448822 -4186
rect 448266 -4742 448502 -4506
rect 448586 -4742 448822 -4506
rect 441986 -7302 442222 -7066
rect 442306 -7302 442542 -7066
rect 441986 -7622 442222 -7386
rect 442306 -7622 442542 -7386
rect 454546 707482 454782 707718
rect 454866 707482 455102 707718
rect 454546 707162 454782 707398
rect 454866 707162 455102 707398
rect 454546 672938 454782 673174
rect 454866 672938 455102 673174
rect 454546 672618 454782 672854
rect 454866 672618 455102 672854
rect 454546 636938 454782 637174
rect 454866 636938 455102 637174
rect 454546 636618 454782 636854
rect 454866 636618 455102 636854
rect 454546 600938 454782 601174
rect 454866 600938 455102 601174
rect 454546 600618 454782 600854
rect 454866 600618 455102 600854
rect 454546 564938 454782 565174
rect 454866 564938 455102 565174
rect 454546 564618 454782 564854
rect 454866 564618 455102 564854
rect 454546 528938 454782 529174
rect 454866 528938 455102 529174
rect 454546 528618 454782 528854
rect 454866 528618 455102 528854
rect 454546 492938 454782 493174
rect 454866 492938 455102 493174
rect 454546 492618 454782 492854
rect 454866 492618 455102 492854
rect 454546 456938 454782 457174
rect 454866 456938 455102 457174
rect 454546 456618 454782 456854
rect 454866 456618 455102 456854
rect 454546 420938 454782 421174
rect 454866 420938 455102 421174
rect 454546 420618 454782 420854
rect 454866 420618 455102 420854
rect 454546 384938 454782 385174
rect 454866 384938 455102 385174
rect 454546 384618 454782 384854
rect 454866 384618 455102 384854
rect 454546 348938 454782 349174
rect 454866 348938 455102 349174
rect 454546 348618 454782 348854
rect 454866 348618 455102 348854
rect 454546 312938 454782 313174
rect 454866 312938 455102 313174
rect 454546 312618 454782 312854
rect 454866 312618 455102 312854
rect 454546 276938 454782 277174
rect 454866 276938 455102 277174
rect 454546 276618 454782 276854
rect 454866 276618 455102 276854
rect 454546 240938 454782 241174
rect 454866 240938 455102 241174
rect 454546 240618 454782 240854
rect 454866 240618 455102 240854
rect 454546 204938 454782 205174
rect 454866 204938 455102 205174
rect 454546 204618 454782 204854
rect 454866 204618 455102 204854
rect 454546 168938 454782 169174
rect 454866 168938 455102 169174
rect 454546 168618 454782 168854
rect 454866 168618 455102 168854
rect 454546 132938 454782 133174
rect 454866 132938 455102 133174
rect 454546 132618 454782 132854
rect 454866 132618 455102 132854
rect 454546 96938 454782 97174
rect 454866 96938 455102 97174
rect 454546 96618 454782 96854
rect 454866 96618 455102 96854
rect 454546 60938 454782 61174
rect 454866 60938 455102 61174
rect 454546 60618 454782 60854
rect 454866 60618 455102 60854
rect 454546 24938 454782 25174
rect 454866 24938 455102 25174
rect 454546 24618 454782 24854
rect 454866 24618 455102 24854
rect 454546 -3462 454782 -3226
rect 454866 -3462 455102 -3226
rect 454546 -3782 454782 -3546
rect 454866 -3782 455102 -3546
rect 458266 676658 458502 676894
rect 458586 676658 458822 676894
rect 458266 676338 458502 676574
rect 458586 676338 458822 676574
rect 458266 640658 458502 640894
rect 458586 640658 458822 640894
rect 458266 640338 458502 640574
rect 458586 640338 458822 640574
rect 458266 604658 458502 604894
rect 458586 604658 458822 604894
rect 458266 604338 458502 604574
rect 458586 604338 458822 604574
rect 458266 568658 458502 568894
rect 458586 568658 458822 568894
rect 458266 568338 458502 568574
rect 458586 568338 458822 568574
rect 458266 532658 458502 532894
rect 458586 532658 458822 532894
rect 458266 532338 458502 532574
rect 458586 532338 458822 532574
rect 458266 496658 458502 496894
rect 458586 496658 458822 496894
rect 458266 496338 458502 496574
rect 458586 496338 458822 496574
rect 458266 460658 458502 460894
rect 458586 460658 458822 460894
rect 458266 460338 458502 460574
rect 458586 460338 458822 460574
rect 458266 424658 458502 424894
rect 458586 424658 458822 424894
rect 458266 424338 458502 424574
rect 458586 424338 458822 424574
rect 458266 388658 458502 388894
rect 458586 388658 458822 388894
rect 458266 388338 458502 388574
rect 458586 388338 458822 388574
rect 458266 352658 458502 352894
rect 458586 352658 458822 352894
rect 458266 352338 458502 352574
rect 458586 352338 458822 352574
rect 458266 316658 458502 316894
rect 458586 316658 458822 316894
rect 458266 316338 458502 316574
rect 458586 316338 458822 316574
rect 458266 280658 458502 280894
rect 458586 280658 458822 280894
rect 458266 280338 458502 280574
rect 458586 280338 458822 280574
rect 458266 244658 458502 244894
rect 458586 244658 458822 244894
rect 458266 244338 458502 244574
rect 458586 244338 458822 244574
rect 458266 208658 458502 208894
rect 458586 208658 458822 208894
rect 458266 208338 458502 208574
rect 458586 208338 458822 208574
rect 458266 172658 458502 172894
rect 458586 172658 458822 172894
rect 458266 172338 458502 172574
rect 458586 172338 458822 172574
rect 458266 136658 458502 136894
rect 458586 136658 458822 136894
rect 458266 136338 458502 136574
rect 458586 136338 458822 136574
rect 458266 100658 458502 100894
rect 458586 100658 458822 100894
rect 458266 100338 458502 100574
rect 458586 100338 458822 100574
rect 458266 64658 458502 64894
rect 458586 64658 458822 64894
rect 458266 64338 458502 64574
rect 458586 64338 458822 64574
rect 458266 28658 458502 28894
rect 458586 28658 458822 28894
rect 458266 28338 458502 28574
rect 458586 28338 458822 28574
rect 460826 704602 461062 704838
rect 461146 704602 461382 704838
rect 460826 704282 461062 704518
rect 461146 704282 461382 704518
rect 460826 687218 461062 687454
rect 461146 687218 461382 687454
rect 460826 686898 461062 687134
rect 461146 686898 461382 687134
rect 460826 651218 461062 651454
rect 461146 651218 461382 651454
rect 460826 650898 461062 651134
rect 461146 650898 461382 651134
rect 460826 615218 461062 615454
rect 461146 615218 461382 615454
rect 460826 614898 461062 615134
rect 461146 614898 461382 615134
rect 460826 579218 461062 579454
rect 461146 579218 461382 579454
rect 460826 578898 461062 579134
rect 461146 578898 461382 579134
rect 460826 543218 461062 543454
rect 461146 543218 461382 543454
rect 460826 542898 461062 543134
rect 461146 542898 461382 543134
rect 460826 507218 461062 507454
rect 461146 507218 461382 507454
rect 460826 506898 461062 507134
rect 461146 506898 461382 507134
rect 460826 471218 461062 471454
rect 461146 471218 461382 471454
rect 460826 470898 461062 471134
rect 461146 470898 461382 471134
rect 460826 435218 461062 435454
rect 461146 435218 461382 435454
rect 460826 434898 461062 435134
rect 461146 434898 461382 435134
rect 460826 399218 461062 399454
rect 461146 399218 461382 399454
rect 460826 398898 461062 399134
rect 461146 398898 461382 399134
rect 460826 363218 461062 363454
rect 461146 363218 461382 363454
rect 460826 362898 461062 363134
rect 461146 362898 461382 363134
rect 460826 327218 461062 327454
rect 461146 327218 461382 327454
rect 460826 326898 461062 327134
rect 461146 326898 461382 327134
rect 460826 291218 461062 291454
rect 461146 291218 461382 291454
rect 460826 290898 461062 291134
rect 461146 290898 461382 291134
rect 460826 255218 461062 255454
rect 461146 255218 461382 255454
rect 460826 254898 461062 255134
rect 461146 254898 461382 255134
rect 460826 219218 461062 219454
rect 461146 219218 461382 219454
rect 460826 218898 461062 219134
rect 461146 218898 461382 219134
rect 460826 183218 461062 183454
rect 461146 183218 461382 183454
rect 460826 182898 461062 183134
rect 461146 182898 461382 183134
rect 460826 147218 461062 147454
rect 461146 147218 461382 147454
rect 460826 146898 461062 147134
rect 461146 146898 461382 147134
rect 460826 111218 461062 111454
rect 461146 111218 461382 111454
rect 460826 110898 461062 111134
rect 461146 110898 461382 111134
rect 460826 75218 461062 75454
rect 461146 75218 461382 75454
rect 460826 74898 461062 75134
rect 461146 74898 461382 75134
rect 460826 39218 461062 39454
rect 461146 39218 461382 39454
rect 460826 38898 461062 39134
rect 461146 38898 461382 39134
rect 460826 3218 461062 3454
rect 461146 3218 461382 3454
rect 460826 2898 461062 3134
rect 461146 2898 461382 3134
rect 460826 -582 461062 -346
rect 461146 -582 461382 -346
rect 460826 -902 461062 -666
rect 461146 -902 461382 -666
rect 471986 710362 472222 710598
rect 472306 710362 472542 710598
rect 471986 710042 472222 710278
rect 472306 710042 472542 710278
rect 468266 708442 468502 708678
rect 468586 708442 468822 708678
rect 468266 708122 468502 708358
rect 468586 708122 468822 708358
rect 461986 680378 462222 680614
rect 462306 680378 462542 680614
rect 461986 680058 462222 680294
rect 462306 680058 462542 680294
rect 461986 644378 462222 644614
rect 462306 644378 462542 644614
rect 461986 644058 462222 644294
rect 462306 644058 462542 644294
rect 461986 608378 462222 608614
rect 462306 608378 462542 608614
rect 461986 608058 462222 608294
rect 462306 608058 462542 608294
rect 461986 572378 462222 572614
rect 462306 572378 462542 572614
rect 461986 572058 462222 572294
rect 462306 572058 462542 572294
rect 461986 536378 462222 536614
rect 462306 536378 462542 536614
rect 461986 536058 462222 536294
rect 462306 536058 462542 536294
rect 461986 500378 462222 500614
rect 462306 500378 462542 500614
rect 461986 500058 462222 500294
rect 462306 500058 462542 500294
rect 461986 464378 462222 464614
rect 462306 464378 462542 464614
rect 461986 464058 462222 464294
rect 462306 464058 462542 464294
rect 461986 428378 462222 428614
rect 462306 428378 462542 428614
rect 461986 428058 462222 428294
rect 462306 428058 462542 428294
rect 461986 392378 462222 392614
rect 462306 392378 462542 392614
rect 461986 392058 462222 392294
rect 462306 392058 462542 392294
rect 461986 356378 462222 356614
rect 462306 356378 462542 356614
rect 461986 356058 462222 356294
rect 462306 356058 462542 356294
rect 461986 320378 462222 320614
rect 462306 320378 462542 320614
rect 461986 320058 462222 320294
rect 462306 320058 462542 320294
rect 461986 284378 462222 284614
rect 462306 284378 462542 284614
rect 461986 284058 462222 284294
rect 462306 284058 462542 284294
rect 461986 248378 462222 248614
rect 462306 248378 462542 248614
rect 461986 248058 462222 248294
rect 462306 248058 462542 248294
rect 461986 212378 462222 212614
rect 462306 212378 462542 212614
rect 461986 212058 462222 212294
rect 462306 212058 462542 212294
rect 461986 176378 462222 176614
rect 462306 176378 462542 176614
rect 461986 176058 462222 176294
rect 462306 176058 462542 176294
rect 461986 140378 462222 140614
rect 462306 140378 462542 140614
rect 461986 140058 462222 140294
rect 462306 140058 462542 140294
rect 461986 104378 462222 104614
rect 462306 104378 462542 104614
rect 461986 104058 462222 104294
rect 462306 104058 462542 104294
rect 461986 68378 462222 68614
rect 462306 68378 462542 68614
rect 461986 68058 462222 68294
rect 462306 68058 462542 68294
rect 461986 32378 462222 32614
rect 462306 32378 462542 32614
rect 461986 32058 462222 32294
rect 462306 32058 462542 32294
rect 458266 -5382 458502 -5146
rect 458586 -5382 458822 -5146
rect 458266 -5702 458502 -5466
rect 458586 -5702 458822 -5466
rect 451986 -6342 452222 -6106
rect 452306 -6342 452542 -6106
rect 451986 -6662 452222 -6426
rect 452306 -6662 452542 -6426
rect 464546 706522 464782 706758
rect 464866 706522 465102 706758
rect 464546 706202 464782 706438
rect 464866 706202 465102 706438
rect 464546 690938 464782 691174
rect 464866 690938 465102 691174
rect 464546 690618 464782 690854
rect 464866 690618 465102 690854
rect 464546 654938 464782 655174
rect 464866 654938 465102 655174
rect 464546 654618 464782 654854
rect 464866 654618 465102 654854
rect 464546 618938 464782 619174
rect 464866 618938 465102 619174
rect 464546 618618 464782 618854
rect 464866 618618 465102 618854
rect 464546 582938 464782 583174
rect 464866 582938 465102 583174
rect 464546 582618 464782 582854
rect 464866 582618 465102 582854
rect 464546 546938 464782 547174
rect 464866 546938 465102 547174
rect 464546 546618 464782 546854
rect 464866 546618 465102 546854
rect 464546 510938 464782 511174
rect 464866 510938 465102 511174
rect 464546 510618 464782 510854
rect 464866 510618 465102 510854
rect 464546 474938 464782 475174
rect 464866 474938 465102 475174
rect 464546 474618 464782 474854
rect 464866 474618 465102 474854
rect 464546 438938 464782 439174
rect 464866 438938 465102 439174
rect 464546 438618 464782 438854
rect 464866 438618 465102 438854
rect 464546 402938 464782 403174
rect 464866 402938 465102 403174
rect 464546 402618 464782 402854
rect 464866 402618 465102 402854
rect 464546 366938 464782 367174
rect 464866 366938 465102 367174
rect 464546 366618 464782 366854
rect 464866 366618 465102 366854
rect 464546 330938 464782 331174
rect 464866 330938 465102 331174
rect 464546 330618 464782 330854
rect 464866 330618 465102 330854
rect 464546 294938 464782 295174
rect 464866 294938 465102 295174
rect 464546 294618 464782 294854
rect 464866 294618 465102 294854
rect 464546 258938 464782 259174
rect 464866 258938 465102 259174
rect 464546 258618 464782 258854
rect 464866 258618 465102 258854
rect 464546 222938 464782 223174
rect 464866 222938 465102 223174
rect 464546 222618 464782 222854
rect 464866 222618 465102 222854
rect 464546 186938 464782 187174
rect 464866 186938 465102 187174
rect 464546 186618 464782 186854
rect 464866 186618 465102 186854
rect 464546 150938 464782 151174
rect 464866 150938 465102 151174
rect 464546 150618 464782 150854
rect 464866 150618 465102 150854
rect 464546 114938 464782 115174
rect 464866 114938 465102 115174
rect 464546 114618 464782 114854
rect 464866 114618 465102 114854
rect 464546 78938 464782 79174
rect 464866 78938 465102 79174
rect 464546 78618 464782 78854
rect 464866 78618 465102 78854
rect 464546 42938 464782 43174
rect 464866 42938 465102 43174
rect 464546 42618 464782 42854
rect 464866 42618 465102 42854
rect 464546 6938 464782 7174
rect 464866 6938 465102 7174
rect 464546 6618 464782 6854
rect 464866 6618 465102 6854
rect 464546 -2502 464782 -2266
rect 464866 -2502 465102 -2266
rect 464546 -2822 464782 -2586
rect 464866 -2822 465102 -2586
rect 468266 694658 468502 694894
rect 468586 694658 468822 694894
rect 468266 694338 468502 694574
rect 468586 694338 468822 694574
rect 468266 658658 468502 658894
rect 468586 658658 468822 658894
rect 468266 658338 468502 658574
rect 468586 658338 468822 658574
rect 468266 622658 468502 622894
rect 468586 622658 468822 622894
rect 468266 622338 468502 622574
rect 468586 622338 468822 622574
rect 468266 586658 468502 586894
rect 468586 586658 468822 586894
rect 468266 586338 468502 586574
rect 468586 586338 468822 586574
rect 468266 550658 468502 550894
rect 468586 550658 468822 550894
rect 468266 550338 468502 550574
rect 468586 550338 468822 550574
rect 468266 514658 468502 514894
rect 468586 514658 468822 514894
rect 468266 514338 468502 514574
rect 468586 514338 468822 514574
rect 468266 478658 468502 478894
rect 468586 478658 468822 478894
rect 468266 478338 468502 478574
rect 468586 478338 468822 478574
rect 468266 442658 468502 442894
rect 468586 442658 468822 442894
rect 468266 442338 468502 442574
rect 468586 442338 468822 442574
rect 468266 406658 468502 406894
rect 468586 406658 468822 406894
rect 468266 406338 468502 406574
rect 468586 406338 468822 406574
rect 468266 370658 468502 370894
rect 468586 370658 468822 370894
rect 468266 370338 468502 370574
rect 468586 370338 468822 370574
rect 468266 334658 468502 334894
rect 468586 334658 468822 334894
rect 468266 334338 468502 334574
rect 468586 334338 468822 334574
rect 468266 298658 468502 298894
rect 468586 298658 468822 298894
rect 468266 298338 468502 298574
rect 468586 298338 468822 298574
rect 468266 262658 468502 262894
rect 468586 262658 468822 262894
rect 468266 262338 468502 262574
rect 468586 262338 468822 262574
rect 468266 226658 468502 226894
rect 468586 226658 468822 226894
rect 468266 226338 468502 226574
rect 468586 226338 468822 226574
rect 468266 190658 468502 190894
rect 468586 190658 468822 190894
rect 468266 190338 468502 190574
rect 468586 190338 468822 190574
rect 468266 154658 468502 154894
rect 468586 154658 468822 154894
rect 468266 154338 468502 154574
rect 468586 154338 468822 154574
rect 468266 118658 468502 118894
rect 468586 118658 468822 118894
rect 468266 118338 468502 118574
rect 468586 118338 468822 118574
rect 468266 82658 468502 82894
rect 468586 82658 468822 82894
rect 468266 82338 468502 82574
rect 468586 82338 468822 82574
rect 468266 46658 468502 46894
rect 468586 46658 468822 46894
rect 468266 46338 468502 46574
rect 468586 46338 468822 46574
rect 468266 10658 468502 10894
rect 468586 10658 468822 10894
rect 468266 10338 468502 10574
rect 468586 10338 468822 10574
rect 470826 705562 471062 705798
rect 471146 705562 471382 705798
rect 470826 705242 471062 705478
rect 471146 705242 471382 705478
rect 470826 669218 471062 669454
rect 471146 669218 471382 669454
rect 470826 668898 471062 669134
rect 471146 668898 471382 669134
rect 470826 633218 471062 633454
rect 471146 633218 471382 633454
rect 470826 632898 471062 633134
rect 471146 632898 471382 633134
rect 470826 597218 471062 597454
rect 471146 597218 471382 597454
rect 470826 596898 471062 597134
rect 471146 596898 471382 597134
rect 470826 561218 471062 561454
rect 471146 561218 471382 561454
rect 470826 560898 471062 561134
rect 471146 560898 471382 561134
rect 470826 525218 471062 525454
rect 471146 525218 471382 525454
rect 470826 524898 471062 525134
rect 471146 524898 471382 525134
rect 470826 489218 471062 489454
rect 471146 489218 471382 489454
rect 470826 488898 471062 489134
rect 471146 488898 471382 489134
rect 470826 453218 471062 453454
rect 471146 453218 471382 453454
rect 470826 452898 471062 453134
rect 471146 452898 471382 453134
rect 470826 417218 471062 417454
rect 471146 417218 471382 417454
rect 470826 416898 471062 417134
rect 471146 416898 471382 417134
rect 470826 381218 471062 381454
rect 471146 381218 471382 381454
rect 470826 380898 471062 381134
rect 471146 380898 471382 381134
rect 470826 345218 471062 345454
rect 471146 345218 471382 345454
rect 470826 344898 471062 345134
rect 471146 344898 471382 345134
rect 470826 309218 471062 309454
rect 471146 309218 471382 309454
rect 470826 308898 471062 309134
rect 471146 308898 471382 309134
rect 470826 273218 471062 273454
rect 471146 273218 471382 273454
rect 470826 272898 471062 273134
rect 471146 272898 471382 273134
rect 470826 237218 471062 237454
rect 471146 237218 471382 237454
rect 470826 236898 471062 237134
rect 471146 236898 471382 237134
rect 470826 201218 471062 201454
rect 471146 201218 471382 201454
rect 470826 200898 471062 201134
rect 471146 200898 471382 201134
rect 470826 165218 471062 165454
rect 471146 165218 471382 165454
rect 470826 164898 471062 165134
rect 471146 164898 471382 165134
rect 470826 129218 471062 129454
rect 471146 129218 471382 129454
rect 470826 128898 471062 129134
rect 471146 128898 471382 129134
rect 470826 93218 471062 93454
rect 471146 93218 471382 93454
rect 470826 92898 471062 93134
rect 471146 92898 471382 93134
rect 470826 57218 471062 57454
rect 471146 57218 471382 57454
rect 470826 56898 471062 57134
rect 471146 56898 471382 57134
rect 470826 21218 471062 21454
rect 471146 21218 471382 21454
rect 470826 20898 471062 21134
rect 471146 20898 471382 21134
rect 470826 -1542 471062 -1306
rect 471146 -1542 471382 -1306
rect 470826 -1862 471062 -1626
rect 471146 -1862 471382 -1626
rect 481986 711322 482222 711558
rect 482306 711322 482542 711558
rect 481986 711002 482222 711238
rect 482306 711002 482542 711238
rect 478266 709402 478502 709638
rect 478586 709402 478822 709638
rect 478266 709082 478502 709318
rect 478586 709082 478822 709318
rect 471986 698378 472222 698614
rect 472306 698378 472542 698614
rect 471986 698058 472222 698294
rect 472306 698058 472542 698294
rect 471986 662378 472222 662614
rect 472306 662378 472542 662614
rect 471986 662058 472222 662294
rect 472306 662058 472542 662294
rect 471986 626378 472222 626614
rect 472306 626378 472542 626614
rect 471986 626058 472222 626294
rect 472306 626058 472542 626294
rect 471986 590378 472222 590614
rect 472306 590378 472542 590614
rect 471986 590058 472222 590294
rect 472306 590058 472542 590294
rect 471986 554378 472222 554614
rect 472306 554378 472542 554614
rect 471986 554058 472222 554294
rect 472306 554058 472542 554294
rect 471986 518378 472222 518614
rect 472306 518378 472542 518614
rect 471986 518058 472222 518294
rect 472306 518058 472542 518294
rect 471986 482378 472222 482614
rect 472306 482378 472542 482614
rect 471986 482058 472222 482294
rect 472306 482058 472542 482294
rect 471986 446378 472222 446614
rect 472306 446378 472542 446614
rect 471986 446058 472222 446294
rect 472306 446058 472542 446294
rect 471986 410378 472222 410614
rect 472306 410378 472542 410614
rect 471986 410058 472222 410294
rect 472306 410058 472542 410294
rect 471986 374378 472222 374614
rect 472306 374378 472542 374614
rect 471986 374058 472222 374294
rect 472306 374058 472542 374294
rect 471986 338378 472222 338614
rect 472306 338378 472542 338614
rect 471986 338058 472222 338294
rect 472306 338058 472542 338294
rect 471986 302378 472222 302614
rect 472306 302378 472542 302614
rect 471986 302058 472222 302294
rect 472306 302058 472542 302294
rect 471986 266378 472222 266614
rect 472306 266378 472542 266614
rect 471986 266058 472222 266294
rect 472306 266058 472542 266294
rect 471986 230378 472222 230614
rect 472306 230378 472542 230614
rect 471986 230058 472222 230294
rect 472306 230058 472542 230294
rect 471986 194378 472222 194614
rect 472306 194378 472542 194614
rect 471986 194058 472222 194294
rect 472306 194058 472542 194294
rect 471986 158378 472222 158614
rect 472306 158378 472542 158614
rect 471986 158058 472222 158294
rect 472306 158058 472542 158294
rect 471986 122378 472222 122614
rect 472306 122378 472542 122614
rect 471986 122058 472222 122294
rect 472306 122058 472542 122294
rect 471986 86378 472222 86614
rect 472306 86378 472542 86614
rect 471986 86058 472222 86294
rect 472306 86058 472542 86294
rect 471986 50378 472222 50614
rect 472306 50378 472542 50614
rect 471986 50058 472222 50294
rect 472306 50058 472542 50294
rect 471986 14378 472222 14614
rect 472306 14378 472542 14614
rect 471986 14058 472222 14294
rect 472306 14058 472542 14294
rect 468266 -4422 468502 -4186
rect 468586 -4422 468822 -4186
rect 468266 -4742 468502 -4506
rect 468586 -4742 468822 -4506
rect 461986 -7302 462222 -7066
rect 462306 -7302 462542 -7066
rect 461986 -7622 462222 -7386
rect 462306 -7622 462542 -7386
rect 474546 707482 474782 707718
rect 474866 707482 475102 707718
rect 474546 707162 474782 707398
rect 474866 707162 475102 707398
rect 474546 672938 474782 673174
rect 474866 672938 475102 673174
rect 474546 672618 474782 672854
rect 474866 672618 475102 672854
rect 474546 636938 474782 637174
rect 474866 636938 475102 637174
rect 474546 636618 474782 636854
rect 474866 636618 475102 636854
rect 474546 600938 474782 601174
rect 474866 600938 475102 601174
rect 474546 600618 474782 600854
rect 474866 600618 475102 600854
rect 474546 564938 474782 565174
rect 474866 564938 475102 565174
rect 474546 564618 474782 564854
rect 474866 564618 475102 564854
rect 474546 528938 474782 529174
rect 474866 528938 475102 529174
rect 474546 528618 474782 528854
rect 474866 528618 475102 528854
rect 474546 492938 474782 493174
rect 474866 492938 475102 493174
rect 474546 492618 474782 492854
rect 474866 492618 475102 492854
rect 474546 456938 474782 457174
rect 474866 456938 475102 457174
rect 474546 456618 474782 456854
rect 474866 456618 475102 456854
rect 474546 420938 474782 421174
rect 474866 420938 475102 421174
rect 474546 420618 474782 420854
rect 474866 420618 475102 420854
rect 474546 384938 474782 385174
rect 474866 384938 475102 385174
rect 474546 384618 474782 384854
rect 474866 384618 475102 384854
rect 474546 348938 474782 349174
rect 474866 348938 475102 349174
rect 474546 348618 474782 348854
rect 474866 348618 475102 348854
rect 474546 312938 474782 313174
rect 474866 312938 475102 313174
rect 474546 312618 474782 312854
rect 474866 312618 475102 312854
rect 474546 276938 474782 277174
rect 474866 276938 475102 277174
rect 474546 276618 474782 276854
rect 474866 276618 475102 276854
rect 474546 240938 474782 241174
rect 474866 240938 475102 241174
rect 474546 240618 474782 240854
rect 474866 240618 475102 240854
rect 474546 204938 474782 205174
rect 474866 204938 475102 205174
rect 474546 204618 474782 204854
rect 474866 204618 475102 204854
rect 474546 168938 474782 169174
rect 474866 168938 475102 169174
rect 474546 168618 474782 168854
rect 474866 168618 475102 168854
rect 474546 132938 474782 133174
rect 474866 132938 475102 133174
rect 474546 132618 474782 132854
rect 474866 132618 475102 132854
rect 474546 96938 474782 97174
rect 474866 96938 475102 97174
rect 474546 96618 474782 96854
rect 474866 96618 475102 96854
rect 474546 60938 474782 61174
rect 474866 60938 475102 61174
rect 474546 60618 474782 60854
rect 474866 60618 475102 60854
rect 474546 24938 474782 25174
rect 474866 24938 475102 25174
rect 474546 24618 474782 24854
rect 474866 24618 475102 24854
rect 474546 -3462 474782 -3226
rect 474866 -3462 475102 -3226
rect 474546 -3782 474782 -3546
rect 474866 -3782 475102 -3546
rect 478266 676658 478502 676894
rect 478586 676658 478822 676894
rect 478266 676338 478502 676574
rect 478586 676338 478822 676574
rect 478266 640658 478502 640894
rect 478586 640658 478822 640894
rect 478266 640338 478502 640574
rect 478586 640338 478822 640574
rect 478266 604658 478502 604894
rect 478586 604658 478822 604894
rect 478266 604338 478502 604574
rect 478586 604338 478822 604574
rect 478266 568658 478502 568894
rect 478586 568658 478822 568894
rect 478266 568338 478502 568574
rect 478586 568338 478822 568574
rect 478266 532658 478502 532894
rect 478586 532658 478822 532894
rect 478266 532338 478502 532574
rect 478586 532338 478822 532574
rect 478266 496658 478502 496894
rect 478586 496658 478822 496894
rect 478266 496338 478502 496574
rect 478586 496338 478822 496574
rect 478266 460658 478502 460894
rect 478586 460658 478822 460894
rect 478266 460338 478502 460574
rect 478586 460338 478822 460574
rect 478266 424658 478502 424894
rect 478586 424658 478822 424894
rect 478266 424338 478502 424574
rect 478586 424338 478822 424574
rect 478266 388658 478502 388894
rect 478586 388658 478822 388894
rect 478266 388338 478502 388574
rect 478586 388338 478822 388574
rect 478266 352658 478502 352894
rect 478586 352658 478822 352894
rect 478266 352338 478502 352574
rect 478586 352338 478822 352574
rect 478266 316658 478502 316894
rect 478586 316658 478822 316894
rect 478266 316338 478502 316574
rect 478586 316338 478822 316574
rect 478266 280658 478502 280894
rect 478586 280658 478822 280894
rect 478266 280338 478502 280574
rect 478586 280338 478822 280574
rect 478266 244658 478502 244894
rect 478586 244658 478822 244894
rect 478266 244338 478502 244574
rect 478586 244338 478822 244574
rect 478266 208658 478502 208894
rect 478586 208658 478822 208894
rect 478266 208338 478502 208574
rect 478586 208338 478822 208574
rect 478266 172658 478502 172894
rect 478586 172658 478822 172894
rect 478266 172338 478502 172574
rect 478586 172338 478822 172574
rect 478266 136658 478502 136894
rect 478586 136658 478822 136894
rect 478266 136338 478502 136574
rect 478586 136338 478822 136574
rect 478266 100658 478502 100894
rect 478586 100658 478822 100894
rect 478266 100338 478502 100574
rect 478586 100338 478822 100574
rect 478266 64658 478502 64894
rect 478586 64658 478822 64894
rect 478266 64338 478502 64574
rect 478586 64338 478822 64574
rect 478266 28658 478502 28894
rect 478586 28658 478822 28894
rect 478266 28338 478502 28574
rect 478586 28338 478822 28574
rect 480826 704602 481062 704838
rect 481146 704602 481382 704838
rect 480826 704282 481062 704518
rect 481146 704282 481382 704518
rect 480826 687218 481062 687454
rect 481146 687218 481382 687454
rect 480826 686898 481062 687134
rect 481146 686898 481382 687134
rect 480826 651218 481062 651454
rect 481146 651218 481382 651454
rect 480826 650898 481062 651134
rect 481146 650898 481382 651134
rect 480826 615218 481062 615454
rect 481146 615218 481382 615454
rect 480826 614898 481062 615134
rect 481146 614898 481382 615134
rect 480826 579218 481062 579454
rect 481146 579218 481382 579454
rect 480826 578898 481062 579134
rect 481146 578898 481382 579134
rect 480826 543218 481062 543454
rect 481146 543218 481382 543454
rect 480826 542898 481062 543134
rect 481146 542898 481382 543134
rect 480826 507218 481062 507454
rect 481146 507218 481382 507454
rect 480826 506898 481062 507134
rect 481146 506898 481382 507134
rect 480826 471218 481062 471454
rect 481146 471218 481382 471454
rect 480826 470898 481062 471134
rect 481146 470898 481382 471134
rect 480826 435218 481062 435454
rect 481146 435218 481382 435454
rect 480826 434898 481062 435134
rect 481146 434898 481382 435134
rect 480826 399218 481062 399454
rect 481146 399218 481382 399454
rect 480826 398898 481062 399134
rect 481146 398898 481382 399134
rect 480826 363218 481062 363454
rect 481146 363218 481382 363454
rect 480826 362898 481062 363134
rect 481146 362898 481382 363134
rect 480826 327218 481062 327454
rect 481146 327218 481382 327454
rect 480826 326898 481062 327134
rect 481146 326898 481382 327134
rect 480826 291218 481062 291454
rect 481146 291218 481382 291454
rect 480826 290898 481062 291134
rect 481146 290898 481382 291134
rect 480826 255218 481062 255454
rect 481146 255218 481382 255454
rect 480826 254898 481062 255134
rect 481146 254898 481382 255134
rect 480826 219218 481062 219454
rect 481146 219218 481382 219454
rect 480826 218898 481062 219134
rect 481146 218898 481382 219134
rect 480826 183218 481062 183454
rect 481146 183218 481382 183454
rect 480826 182898 481062 183134
rect 481146 182898 481382 183134
rect 480826 147218 481062 147454
rect 481146 147218 481382 147454
rect 480826 146898 481062 147134
rect 481146 146898 481382 147134
rect 480826 111218 481062 111454
rect 481146 111218 481382 111454
rect 480826 110898 481062 111134
rect 481146 110898 481382 111134
rect 480826 75218 481062 75454
rect 481146 75218 481382 75454
rect 480826 74898 481062 75134
rect 481146 74898 481382 75134
rect 480826 39218 481062 39454
rect 481146 39218 481382 39454
rect 480826 38898 481062 39134
rect 481146 38898 481382 39134
rect 480826 3218 481062 3454
rect 481146 3218 481382 3454
rect 480826 2898 481062 3134
rect 481146 2898 481382 3134
rect 480826 -582 481062 -346
rect 481146 -582 481382 -346
rect 480826 -902 481062 -666
rect 481146 -902 481382 -666
rect 491986 710362 492222 710598
rect 492306 710362 492542 710598
rect 491986 710042 492222 710278
rect 492306 710042 492542 710278
rect 488266 708442 488502 708678
rect 488586 708442 488822 708678
rect 488266 708122 488502 708358
rect 488586 708122 488822 708358
rect 481986 680378 482222 680614
rect 482306 680378 482542 680614
rect 481986 680058 482222 680294
rect 482306 680058 482542 680294
rect 481986 644378 482222 644614
rect 482306 644378 482542 644614
rect 481986 644058 482222 644294
rect 482306 644058 482542 644294
rect 481986 608378 482222 608614
rect 482306 608378 482542 608614
rect 481986 608058 482222 608294
rect 482306 608058 482542 608294
rect 481986 572378 482222 572614
rect 482306 572378 482542 572614
rect 481986 572058 482222 572294
rect 482306 572058 482542 572294
rect 481986 536378 482222 536614
rect 482306 536378 482542 536614
rect 481986 536058 482222 536294
rect 482306 536058 482542 536294
rect 481986 500378 482222 500614
rect 482306 500378 482542 500614
rect 481986 500058 482222 500294
rect 482306 500058 482542 500294
rect 481986 464378 482222 464614
rect 482306 464378 482542 464614
rect 481986 464058 482222 464294
rect 482306 464058 482542 464294
rect 481986 428378 482222 428614
rect 482306 428378 482542 428614
rect 481986 428058 482222 428294
rect 482306 428058 482542 428294
rect 481986 392378 482222 392614
rect 482306 392378 482542 392614
rect 481986 392058 482222 392294
rect 482306 392058 482542 392294
rect 481986 356378 482222 356614
rect 482306 356378 482542 356614
rect 481986 356058 482222 356294
rect 482306 356058 482542 356294
rect 481986 320378 482222 320614
rect 482306 320378 482542 320614
rect 481986 320058 482222 320294
rect 482306 320058 482542 320294
rect 481986 284378 482222 284614
rect 482306 284378 482542 284614
rect 481986 284058 482222 284294
rect 482306 284058 482542 284294
rect 481986 248378 482222 248614
rect 482306 248378 482542 248614
rect 481986 248058 482222 248294
rect 482306 248058 482542 248294
rect 481986 212378 482222 212614
rect 482306 212378 482542 212614
rect 481986 212058 482222 212294
rect 482306 212058 482542 212294
rect 481986 176378 482222 176614
rect 482306 176378 482542 176614
rect 481986 176058 482222 176294
rect 482306 176058 482542 176294
rect 481986 140378 482222 140614
rect 482306 140378 482542 140614
rect 481986 140058 482222 140294
rect 482306 140058 482542 140294
rect 481986 104378 482222 104614
rect 482306 104378 482542 104614
rect 481986 104058 482222 104294
rect 482306 104058 482542 104294
rect 481986 68378 482222 68614
rect 482306 68378 482542 68614
rect 481986 68058 482222 68294
rect 482306 68058 482542 68294
rect 481986 32378 482222 32614
rect 482306 32378 482542 32614
rect 481986 32058 482222 32294
rect 482306 32058 482542 32294
rect 478266 -5382 478502 -5146
rect 478586 -5382 478822 -5146
rect 478266 -5702 478502 -5466
rect 478586 -5702 478822 -5466
rect 471986 -6342 472222 -6106
rect 472306 -6342 472542 -6106
rect 471986 -6662 472222 -6426
rect 472306 -6662 472542 -6426
rect 484546 706522 484782 706758
rect 484866 706522 485102 706758
rect 484546 706202 484782 706438
rect 484866 706202 485102 706438
rect 484546 690938 484782 691174
rect 484866 690938 485102 691174
rect 484546 690618 484782 690854
rect 484866 690618 485102 690854
rect 484546 654938 484782 655174
rect 484866 654938 485102 655174
rect 484546 654618 484782 654854
rect 484866 654618 485102 654854
rect 484546 618938 484782 619174
rect 484866 618938 485102 619174
rect 484546 618618 484782 618854
rect 484866 618618 485102 618854
rect 484546 582938 484782 583174
rect 484866 582938 485102 583174
rect 484546 582618 484782 582854
rect 484866 582618 485102 582854
rect 484546 546938 484782 547174
rect 484866 546938 485102 547174
rect 484546 546618 484782 546854
rect 484866 546618 485102 546854
rect 484546 510938 484782 511174
rect 484866 510938 485102 511174
rect 484546 510618 484782 510854
rect 484866 510618 485102 510854
rect 484546 474938 484782 475174
rect 484866 474938 485102 475174
rect 484546 474618 484782 474854
rect 484866 474618 485102 474854
rect 484546 438938 484782 439174
rect 484866 438938 485102 439174
rect 484546 438618 484782 438854
rect 484866 438618 485102 438854
rect 484546 402938 484782 403174
rect 484866 402938 485102 403174
rect 484546 402618 484782 402854
rect 484866 402618 485102 402854
rect 484546 366938 484782 367174
rect 484866 366938 485102 367174
rect 484546 366618 484782 366854
rect 484866 366618 485102 366854
rect 484546 330938 484782 331174
rect 484866 330938 485102 331174
rect 484546 330618 484782 330854
rect 484866 330618 485102 330854
rect 484546 294938 484782 295174
rect 484866 294938 485102 295174
rect 484546 294618 484782 294854
rect 484866 294618 485102 294854
rect 484546 258938 484782 259174
rect 484866 258938 485102 259174
rect 484546 258618 484782 258854
rect 484866 258618 485102 258854
rect 484546 222938 484782 223174
rect 484866 222938 485102 223174
rect 484546 222618 484782 222854
rect 484866 222618 485102 222854
rect 484546 186938 484782 187174
rect 484866 186938 485102 187174
rect 484546 186618 484782 186854
rect 484866 186618 485102 186854
rect 484546 150938 484782 151174
rect 484866 150938 485102 151174
rect 484546 150618 484782 150854
rect 484866 150618 485102 150854
rect 484546 114938 484782 115174
rect 484866 114938 485102 115174
rect 484546 114618 484782 114854
rect 484866 114618 485102 114854
rect 484546 78938 484782 79174
rect 484866 78938 485102 79174
rect 484546 78618 484782 78854
rect 484866 78618 485102 78854
rect 484546 42938 484782 43174
rect 484866 42938 485102 43174
rect 484546 42618 484782 42854
rect 484866 42618 485102 42854
rect 484546 6938 484782 7174
rect 484866 6938 485102 7174
rect 484546 6618 484782 6854
rect 484866 6618 485102 6854
rect 484546 -2502 484782 -2266
rect 484866 -2502 485102 -2266
rect 484546 -2822 484782 -2586
rect 484866 -2822 485102 -2586
rect 488266 694658 488502 694894
rect 488586 694658 488822 694894
rect 488266 694338 488502 694574
rect 488586 694338 488822 694574
rect 488266 658658 488502 658894
rect 488586 658658 488822 658894
rect 488266 658338 488502 658574
rect 488586 658338 488822 658574
rect 488266 622658 488502 622894
rect 488586 622658 488822 622894
rect 488266 622338 488502 622574
rect 488586 622338 488822 622574
rect 488266 586658 488502 586894
rect 488586 586658 488822 586894
rect 488266 586338 488502 586574
rect 488586 586338 488822 586574
rect 488266 550658 488502 550894
rect 488586 550658 488822 550894
rect 488266 550338 488502 550574
rect 488586 550338 488822 550574
rect 488266 514658 488502 514894
rect 488586 514658 488822 514894
rect 488266 514338 488502 514574
rect 488586 514338 488822 514574
rect 488266 478658 488502 478894
rect 488586 478658 488822 478894
rect 488266 478338 488502 478574
rect 488586 478338 488822 478574
rect 488266 442658 488502 442894
rect 488586 442658 488822 442894
rect 488266 442338 488502 442574
rect 488586 442338 488822 442574
rect 488266 406658 488502 406894
rect 488586 406658 488822 406894
rect 488266 406338 488502 406574
rect 488586 406338 488822 406574
rect 488266 370658 488502 370894
rect 488586 370658 488822 370894
rect 488266 370338 488502 370574
rect 488586 370338 488822 370574
rect 488266 334658 488502 334894
rect 488586 334658 488822 334894
rect 488266 334338 488502 334574
rect 488586 334338 488822 334574
rect 488266 298658 488502 298894
rect 488586 298658 488822 298894
rect 488266 298338 488502 298574
rect 488586 298338 488822 298574
rect 488266 262658 488502 262894
rect 488586 262658 488822 262894
rect 488266 262338 488502 262574
rect 488586 262338 488822 262574
rect 488266 226658 488502 226894
rect 488586 226658 488822 226894
rect 488266 226338 488502 226574
rect 488586 226338 488822 226574
rect 488266 190658 488502 190894
rect 488586 190658 488822 190894
rect 488266 190338 488502 190574
rect 488586 190338 488822 190574
rect 488266 154658 488502 154894
rect 488586 154658 488822 154894
rect 488266 154338 488502 154574
rect 488586 154338 488822 154574
rect 488266 118658 488502 118894
rect 488586 118658 488822 118894
rect 488266 118338 488502 118574
rect 488586 118338 488822 118574
rect 488266 82658 488502 82894
rect 488586 82658 488822 82894
rect 488266 82338 488502 82574
rect 488586 82338 488822 82574
rect 488266 46658 488502 46894
rect 488586 46658 488822 46894
rect 488266 46338 488502 46574
rect 488586 46338 488822 46574
rect 488266 10658 488502 10894
rect 488586 10658 488822 10894
rect 488266 10338 488502 10574
rect 488586 10338 488822 10574
rect 490826 705562 491062 705798
rect 491146 705562 491382 705798
rect 490826 705242 491062 705478
rect 491146 705242 491382 705478
rect 490826 669218 491062 669454
rect 491146 669218 491382 669454
rect 490826 668898 491062 669134
rect 491146 668898 491382 669134
rect 490826 633218 491062 633454
rect 491146 633218 491382 633454
rect 490826 632898 491062 633134
rect 491146 632898 491382 633134
rect 490826 597218 491062 597454
rect 491146 597218 491382 597454
rect 490826 596898 491062 597134
rect 491146 596898 491382 597134
rect 490826 561218 491062 561454
rect 491146 561218 491382 561454
rect 490826 560898 491062 561134
rect 491146 560898 491382 561134
rect 490826 525218 491062 525454
rect 491146 525218 491382 525454
rect 490826 524898 491062 525134
rect 491146 524898 491382 525134
rect 490826 489218 491062 489454
rect 491146 489218 491382 489454
rect 490826 488898 491062 489134
rect 491146 488898 491382 489134
rect 490826 453218 491062 453454
rect 491146 453218 491382 453454
rect 490826 452898 491062 453134
rect 491146 452898 491382 453134
rect 490826 417218 491062 417454
rect 491146 417218 491382 417454
rect 490826 416898 491062 417134
rect 491146 416898 491382 417134
rect 490826 381218 491062 381454
rect 491146 381218 491382 381454
rect 490826 380898 491062 381134
rect 491146 380898 491382 381134
rect 490826 345218 491062 345454
rect 491146 345218 491382 345454
rect 490826 344898 491062 345134
rect 491146 344898 491382 345134
rect 490826 309218 491062 309454
rect 491146 309218 491382 309454
rect 490826 308898 491062 309134
rect 491146 308898 491382 309134
rect 490826 273218 491062 273454
rect 491146 273218 491382 273454
rect 490826 272898 491062 273134
rect 491146 272898 491382 273134
rect 490826 237218 491062 237454
rect 491146 237218 491382 237454
rect 490826 236898 491062 237134
rect 491146 236898 491382 237134
rect 490826 201218 491062 201454
rect 491146 201218 491382 201454
rect 490826 200898 491062 201134
rect 491146 200898 491382 201134
rect 490826 165218 491062 165454
rect 491146 165218 491382 165454
rect 490826 164898 491062 165134
rect 491146 164898 491382 165134
rect 490826 129218 491062 129454
rect 491146 129218 491382 129454
rect 490826 128898 491062 129134
rect 491146 128898 491382 129134
rect 490826 93218 491062 93454
rect 491146 93218 491382 93454
rect 490826 92898 491062 93134
rect 491146 92898 491382 93134
rect 490826 57218 491062 57454
rect 491146 57218 491382 57454
rect 490826 56898 491062 57134
rect 491146 56898 491382 57134
rect 490826 21218 491062 21454
rect 491146 21218 491382 21454
rect 490826 20898 491062 21134
rect 491146 20898 491382 21134
rect 490826 -1542 491062 -1306
rect 491146 -1542 491382 -1306
rect 490826 -1862 491062 -1626
rect 491146 -1862 491382 -1626
rect 501986 711322 502222 711558
rect 502306 711322 502542 711558
rect 501986 711002 502222 711238
rect 502306 711002 502542 711238
rect 498266 709402 498502 709638
rect 498586 709402 498822 709638
rect 498266 709082 498502 709318
rect 498586 709082 498822 709318
rect 491986 698378 492222 698614
rect 492306 698378 492542 698614
rect 491986 698058 492222 698294
rect 492306 698058 492542 698294
rect 491986 662378 492222 662614
rect 492306 662378 492542 662614
rect 491986 662058 492222 662294
rect 492306 662058 492542 662294
rect 491986 626378 492222 626614
rect 492306 626378 492542 626614
rect 491986 626058 492222 626294
rect 492306 626058 492542 626294
rect 491986 590378 492222 590614
rect 492306 590378 492542 590614
rect 491986 590058 492222 590294
rect 492306 590058 492542 590294
rect 491986 554378 492222 554614
rect 492306 554378 492542 554614
rect 491986 554058 492222 554294
rect 492306 554058 492542 554294
rect 491986 518378 492222 518614
rect 492306 518378 492542 518614
rect 491986 518058 492222 518294
rect 492306 518058 492542 518294
rect 491986 482378 492222 482614
rect 492306 482378 492542 482614
rect 491986 482058 492222 482294
rect 492306 482058 492542 482294
rect 491986 446378 492222 446614
rect 492306 446378 492542 446614
rect 491986 446058 492222 446294
rect 492306 446058 492542 446294
rect 491986 410378 492222 410614
rect 492306 410378 492542 410614
rect 491986 410058 492222 410294
rect 492306 410058 492542 410294
rect 491986 374378 492222 374614
rect 492306 374378 492542 374614
rect 491986 374058 492222 374294
rect 492306 374058 492542 374294
rect 491986 338378 492222 338614
rect 492306 338378 492542 338614
rect 491986 338058 492222 338294
rect 492306 338058 492542 338294
rect 491986 302378 492222 302614
rect 492306 302378 492542 302614
rect 491986 302058 492222 302294
rect 492306 302058 492542 302294
rect 491986 266378 492222 266614
rect 492306 266378 492542 266614
rect 491986 266058 492222 266294
rect 492306 266058 492542 266294
rect 491986 230378 492222 230614
rect 492306 230378 492542 230614
rect 491986 230058 492222 230294
rect 492306 230058 492542 230294
rect 491986 194378 492222 194614
rect 492306 194378 492542 194614
rect 491986 194058 492222 194294
rect 492306 194058 492542 194294
rect 491986 158378 492222 158614
rect 492306 158378 492542 158614
rect 491986 158058 492222 158294
rect 492306 158058 492542 158294
rect 491986 122378 492222 122614
rect 492306 122378 492542 122614
rect 491986 122058 492222 122294
rect 492306 122058 492542 122294
rect 491986 86378 492222 86614
rect 492306 86378 492542 86614
rect 491986 86058 492222 86294
rect 492306 86058 492542 86294
rect 491986 50378 492222 50614
rect 492306 50378 492542 50614
rect 491986 50058 492222 50294
rect 492306 50058 492542 50294
rect 491986 14378 492222 14614
rect 492306 14378 492542 14614
rect 491986 14058 492222 14294
rect 492306 14058 492542 14294
rect 488266 -4422 488502 -4186
rect 488586 -4422 488822 -4186
rect 488266 -4742 488502 -4506
rect 488586 -4742 488822 -4506
rect 481986 -7302 482222 -7066
rect 482306 -7302 482542 -7066
rect 481986 -7622 482222 -7386
rect 482306 -7622 482542 -7386
rect 494546 707482 494782 707718
rect 494866 707482 495102 707718
rect 494546 707162 494782 707398
rect 494866 707162 495102 707398
rect 494546 672938 494782 673174
rect 494866 672938 495102 673174
rect 494546 672618 494782 672854
rect 494866 672618 495102 672854
rect 494546 636938 494782 637174
rect 494866 636938 495102 637174
rect 494546 636618 494782 636854
rect 494866 636618 495102 636854
rect 494546 600938 494782 601174
rect 494866 600938 495102 601174
rect 494546 600618 494782 600854
rect 494866 600618 495102 600854
rect 494546 564938 494782 565174
rect 494866 564938 495102 565174
rect 494546 564618 494782 564854
rect 494866 564618 495102 564854
rect 494546 528938 494782 529174
rect 494866 528938 495102 529174
rect 494546 528618 494782 528854
rect 494866 528618 495102 528854
rect 494546 492938 494782 493174
rect 494866 492938 495102 493174
rect 494546 492618 494782 492854
rect 494866 492618 495102 492854
rect 494546 456938 494782 457174
rect 494866 456938 495102 457174
rect 494546 456618 494782 456854
rect 494866 456618 495102 456854
rect 494546 420938 494782 421174
rect 494866 420938 495102 421174
rect 494546 420618 494782 420854
rect 494866 420618 495102 420854
rect 494546 384938 494782 385174
rect 494866 384938 495102 385174
rect 494546 384618 494782 384854
rect 494866 384618 495102 384854
rect 494546 348938 494782 349174
rect 494866 348938 495102 349174
rect 494546 348618 494782 348854
rect 494866 348618 495102 348854
rect 494546 312938 494782 313174
rect 494866 312938 495102 313174
rect 494546 312618 494782 312854
rect 494866 312618 495102 312854
rect 494546 276938 494782 277174
rect 494866 276938 495102 277174
rect 494546 276618 494782 276854
rect 494866 276618 495102 276854
rect 494546 240938 494782 241174
rect 494866 240938 495102 241174
rect 494546 240618 494782 240854
rect 494866 240618 495102 240854
rect 494546 204938 494782 205174
rect 494866 204938 495102 205174
rect 494546 204618 494782 204854
rect 494866 204618 495102 204854
rect 494546 168938 494782 169174
rect 494866 168938 495102 169174
rect 494546 168618 494782 168854
rect 494866 168618 495102 168854
rect 494546 132938 494782 133174
rect 494866 132938 495102 133174
rect 494546 132618 494782 132854
rect 494866 132618 495102 132854
rect 494546 96938 494782 97174
rect 494866 96938 495102 97174
rect 494546 96618 494782 96854
rect 494866 96618 495102 96854
rect 494546 60938 494782 61174
rect 494866 60938 495102 61174
rect 494546 60618 494782 60854
rect 494866 60618 495102 60854
rect 494546 24938 494782 25174
rect 494866 24938 495102 25174
rect 494546 24618 494782 24854
rect 494866 24618 495102 24854
rect 494546 -3462 494782 -3226
rect 494866 -3462 495102 -3226
rect 494546 -3782 494782 -3546
rect 494866 -3782 495102 -3546
rect 498266 676658 498502 676894
rect 498586 676658 498822 676894
rect 498266 676338 498502 676574
rect 498586 676338 498822 676574
rect 498266 640658 498502 640894
rect 498586 640658 498822 640894
rect 498266 640338 498502 640574
rect 498586 640338 498822 640574
rect 498266 604658 498502 604894
rect 498586 604658 498822 604894
rect 498266 604338 498502 604574
rect 498586 604338 498822 604574
rect 498266 568658 498502 568894
rect 498586 568658 498822 568894
rect 498266 568338 498502 568574
rect 498586 568338 498822 568574
rect 498266 532658 498502 532894
rect 498586 532658 498822 532894
rect 498266 532338 498502 532574
rect 498586 532338 498822 532574
rect 498266 496658 498502 496894
rect 498586 496658 498822 496894
rect 498266 496338 498502 496574
rect 498586 496338 498822 496574
rect 498266 460658 498502 460894
rect 498586 460658 498822 460894
rect 498266 460338 498502 460574
rect 498586 460338 498822 460574
rect 498266 424658 498502 424894
rect 498586 424658 498822 424894
rect 498266 424338 498502 424574
rect 498586 424338 498822 424574
rect 498266 388658 498502 388894
rect 498586 388658 498822 388894
rect 498266 388338 498502 388574
rect 498586 388338 498822 388574
rect 498266 352658 498502 352894
rect 498586 352658 498822 352894
rect 498266 352338 498502 352574
rect 498586 352338 498822 352574
rect 498266 316658 498502 316894
rect 498586 316658 498822 316894
rect 498266 316338 498502 316574
rect 498586 316338 498822 316574
rect 498266 280658 498502 280894
rect 498586 280658 498822 280894
rect 498266 280338 498502 280574
rect 498586 280338 498822 280574
rect 498266 244658 498502 244894
rect 498586 244658 498822 244894
rect 498266 244338 498502 244574
rect 498586 244338 498822 244574
rect 498266 208658 498502 208894
rect 498586 208658 498822 208894
rect 498266 208338 498502 208574
rect 498586 208338 498822 208574
rect 498266 172658 498502 172894
rect 498586 172658 498822 172894
rect 498266 172338 498502 172574
rect 498586 172338 498822 172574
rect 498266 136658 498502 136894
rect 498586 136658 498822 136894
rect 498266 136338 498502 136574
rect 498586 136338 498822 136574
rect 498266 100658 498502 100894
rect 498586 100658 498822 100894
rect 498266 100338 498502 100574
rect 498586 100338 498822 100574
rect 498266 64658 498502 64894
rect 498586 64658 498822 64894
rect 498266 64338 498502 64574
rect 498586 64338 498822 64574
rect 498266 28658 498502 28894
rect 498586 28658 498822 28894
rect 498266 28338 498502 28574
rect 498586 28338 498822 28574
rect 500826 704602 501062 704838
rect 501146 704602 501382 704838
rect 500826 704282 501062 704518
rect 501146 704282 501382 704518
rect 500826 687218 501062 687454
rect 501146 687218 501382 687454
rect 500826 686898 501062 687134
rect 501146 686898 501382 687134
rect 500826 651218 501062 651454
rect 501146 651218 501382 651454
rect 500826 650898 501062 651134
rect 501146 650898 501382 651134
rect 500826 615218 501062 615454
rect 501146 615218 501382 615454
rect 500826 614898 501062 615134
rect 501146 614898 501382 615134
rect 500826 579218 501062 579454
rect 501146 579218 501382 579454
rect 500826 578898 501062 579134
rect 501146 578898 501382 579134
rect 500826 543218 501062 543454
rect 501146 543218 501382 543454
rect 500826 542898 501062 543134
rect 501146 542898 501382 543134
rect 500826 507218 501062 507454
rect 501146 507218 501382 507454
rect 500826 506898 501062 507134
rect 501146 506898 501382 507134
rect 500826 471218 501062 471454
rect 501146 471218 501382 471454
rect 500826 470898 501062 471134
rect 501146 470898 501382 471134
rect 500826 435218 501062 435454
rect 501146 435218 501382 435454
rect 500826 434898 501062 435134
rect 501146 434898 501382 435134
rect 500826 399218 501062 399454
rect 501146 399218 501382 399454
rect 500826 398898 501062 399134
rect 501146 398898 501382 399134
rect 500826 363218 501062 363454
rect 501146 363218 501382 363454
rect 500826 362898 501062 363134
rect 501146 362898 501382 363134
rect 500826 327218 501062 327454
rect 501146 327218 501382 327454
rect 500826 326898 501062 327134
rect 501146 326898 501382 327134
rect 500826 291218 501062 291454
rect 501146 291218 501382 291454
rect 500826 290898 501062 291134
rect 501146 290898 501382 291134
rect 500826 255218 501062 255454
rect 501146 255218 501382 255454
rect 500826 254898 501062 255134
rect 501146 254898 501382 255134
rect 500826 219218 501062 219454
rect 501146 219218 501382 219454
rect 500826 218898 501062 219134
rect 501146 218898 501382 219134
rect 500826 183218 501062 183454
rect 501146 183218 501382 183454
rect 500826 182898 501062 183134
rect 501146 182898 501382 183134
rect 500826 147218 501062 147454
rect 501146 147218 501382 147454
rect 500826 146898 501062 147134
rect 501146 146898 501382 147134
rect 500826 111218 501062 111454
rect 501146 111218 501382 111454
rect 500826 110898 501062 111134
rect 501146 110898 501382 111134
rect 500826 75218 501062 75454
rect 501146 75218 501382 75454
rect 500826 74898 501062 75134
rect 501146 74898 501382 75134
rect 500826 39218 501062 39454
rect 501146 39218 501382 39454
rect 500826 38898 501062 39134
rect 501146 38898 501382 39134
rect 500826 3218 501062 3454
rect 501146 3218 501382 3454
rect 500826 2898 501062 3134
rect 501146 2898 501382 3134
rect 500826 -582 501062 -346
rect 501146 -582 501382 -346
rect 500826 -902 501062 -666
rect 501146 -902 501382 -666
rect 511986 710362 512222 710598
rect 512306 710362 512542 710598
rect 511986 710042 512222 710278
rect 512306 710042 512542 710278
rect 508266 708442 508502 708678
rect 508586 708442 508822 708678
rect 508266 708122 508502 708358
rect 508586 708122 508822 708358
rect 501986 680378 502222 680614
rect 502306 680378 502542 680614
rect 501986 680058 502222 680294
rect 502306 680058 502542 680294
rect 501986 644378 502222 644614
rect 502306 644378 502542 644614
rect 501986 644058 502222 644294
rect 502306 644058 502542 644294
rect 501986 608378 502222 608614
rect 502306 608378 502542 608614
rect 501986 608058 502222 608294
rect 502306 608058 502542 608294
rect 501986 572378 502222 572614
rect 502306 572378 502542 572614
rect 501986 572058 502222 572294
rect 502306 572058 502542 572294
rect 501986 536378 502222 536614
rect 502306 536378 502542 536614
rect 501986 536058 502222 536294
rect 502306 536058 502542 536294
rect 501986 500378 502222 500614
rect 502306 500378 502542 500614
rect 501986 500058 502222 500294
rect 502306 500058 502542 500294
rect 501986 464378 502222 464614
rect 502306 464378 502542 464614
rect 501986 464058 502222 464294
rect 502306 464058 502542 464294
rect 501986 428378 502222 428614
rect 502306 428378 502542 428614
rect 501986 428058 502222 428294
rect 502306 428058 502542 428294
rect 501986 392378 502222 392614
rect 502306 392378 502542 392614
rect 501986 392058 502222 392294
rect 502306 392058 502542 392294
rect 501986 356378 502222 356614
rect 502306 356378 502542 356614
rect 501986 356058 502222 356294
rect 502306 356058 502542 356294
rect 501986 320378 502222 320614
rect 502306 320378 502542 320614
rect 501986 320058 502222 320294
rect 502306 320058 502542 320294
rect 501986 284378 502222 284614
rect 502306 284378 502542 284614
rect 501986 284058 502222 284294
rect 502306 284058 502542 284294
rect 501986 248378 502222 248614
rect 502306 248378 502542 248614
rect 501986 248058 502222 248294
rect 502306 248058 502542 248294
rect 501986 212378 502222 212614
rect 502306 212378 502542 212614
rect 501986 212058 502222 212294
rect 502306 212058 502542 212294
rect 501986 176378 502222 176614
rect 502306 176378 502542 176614
rect 501986 176058 502222 176294
rect 502306 176058 502542 176294
rect 501986 140378 502222 140614
rect 502306 140378 502542 140614
rect 501986 140058 502222 140294
rect 502306 140058 502542 140294
rect 501986 104378 502222 104614
rect 502306 104378 502542 104614
rect 501986 104058 502222 104294
rect 502306 104058 502542 104294
rect 501986 68378 502222 68614
rect 502306 68378 502542 68614
rect 501986 68058 502222 68294
rect 502306 68058 502542 68294
rect 501986 32378 502222 32614
rect 502306 32378 502542 32614
rect 501986 32058 502222 32294
rect 502306 32058 502542 32294
rect 498266 -5382 498502 -5146
rect 498586 -5382 498822 -5146
rect 498266 -5702 498502 -5466
rect 498586 -5702 498822 -5466
rect 491986 -6342 492222 -6106
rect 492306 -6342 492542 -6106
rect 491986 -6662 492222 -6426
rect 492306 -6662 492542 -6426
rect 504546 706522 504782 706758
rect 504866 706522 505102 706758
rect 504546 706202 504782 706438
rect 504866 706202 505102 706438
rect 504546 690938 504782 691174
rect 504866 690938 505102 691174
rect 504546 690618 504782 690854
rect 504866 690618 505102 690854
rect 504546 654938 504782 655174
rect 504866 654938 505102 655174
rect 504546 654618 504782 654854
rect 504866 654618 505102 654854
rect 504546 618938 504782 619174
rect 504866 618938 505102 619174
rect 504546 618618 504782 618854
rect 504866 618618 505102 618854
rect 504546 582938 504782 583174
rect 504866 582938 505102 583174
rect 504546 582618 504782 582854
rect 504866 582618 505102 582854
rect 504546 546938 504782 547174
rect 504866 546938 505102 547174
rect 504546 546618 504782 546854
rect 504866 546618 505102 546854
rect 504546 510938 504782 511174
rect 504866 510938 505102 511174
rect 504546 510618 504782 510854
rect 504866 510618 505102 510854
rect 504546 474938 504782 475174
rect 504866 474938 505102 475174
rect 504546 474618 504782 474854
rect 504866 474618 505102 474854
rect 504546 438938 504782 439174
rect 504866 438938 505102 439174
rect 504546 438618 504782 438854
rect 504866 438618 505102 438854
rect 504546 402938 504782 403174
rect 504866 402938 505102 403174
rect 504546 402618 504782 402854
rect 504866 402618 505102 402854
rect 504546 366938 504782 367174
rect 504866 366938 505102 367174
rect 504546 366618 504782 366854
rect 504866 366618 505102 366854
rect 504546 330938 504782 331174
rect 504866 330938 505102 331174
rect 504546 330618 504782 330854
rect 504866 330618 505102 330854
rect 504546 294938 504782 295174
rect 504866 294938 505102 295174
rect 504546 294618 504782 294854
rect 504866 294618 505102 294854
rect 504546 258938 504782 259174
rect 504866 258938 505102 259174
rect 504546 258618 504782 258854
rect 504866 258618 505102 258854
rect 504546 222938 504782 223174
rect 504866 222938 505102 223174
rect 504546 222618 504782 222854
rect 504866 222618 505102 222854
rect 504546 186938 504782 187174
rect 504866 186938 505102 187174
rect 504546 186618 504782 186854
rect 504866 186618 505102 186854
rect 504546 150938 504782 151174
rect 504866 150938 505102 151174
rect 504546 150618 504782 150854
rect 504866 150618 505102 150854
rect 504546 114938 504782 115174
rect 504866 114938 505102 115174
rect 504546 114618 504782 114854
rect 504866 114618 505102 114854
rect 504546 78938 504782 79174
rect 504866 78938 505102 79174
rect 504546 78618 504782 78854
rect 504866 78618 505102 78854
rect 504546 42938 504782 43174
rect 504866 42938 505102 43174
rect 504546 42618 504782 42854
rect 504866 42618 505102 42854
rect 504546 6938 504782 7174
rect 504866 6938 505102 7174
rect 504546 6618 504782 6854
rect 504866 6618 505102 6854
rect 504546 -2502 504782 -2266
rect 504866 -2502 505102 -2266
rect 504546 -2822 504782 -2586
rect 504866 -2822 505102 -2586
rect 508266 694658 508502 694894
rect 508586 694658 508822 694894
rect 508266 694338 508502 694574
rect 508586 694338 508822 694574
rect 508266 658658 508502 658894
rect 508586 658658 508822 658894
rect 508266 658338 508502 658574
rect 508586 658338 508822 658574
rect 508266 622658 508502 622894
rect 508586 622658 508822 622894
rect 508266 622338 508502 622574
rect 508586 622338 508822 622574
rect 508266 586658 508502 586894
rect 508586 586658 508822 586894
rect 508266 586338 508502 586574
rect 508586 586338 508822 586574
rect 508266 550658 508502 550894
rect 508586 550658 508822 550894
rect 508266 550338 508502 550574
rect 508586 550338 508822 550574
rect 508266 514658 508502 514894
rect 508586 514658 508822 514894
rect 508266 514338 508502 514574
rect 508586 514338 508822 514574
rect 508266 478658 508502 478894
rect 508586 478658 508822 478894
rect 508266 478338 508502 478574
rect 508586 478338 508822 478574
rect 508266 442658 508502 442894
rect 508586 442658 508822 442894
rect 508266 442338 508502 442574
rect 508586 442338 508822 442574
rect 508266 406658 508502 406894
rect 508586 406658 508822 406894
rect 508266 406338 508502 406574
rect 508586 406338 508822 406574
rect 508266 370658 508502 370894
rect 508586 370658 508822 370894
rect 508266 370338 508502 370574
rect 508586 370338 508822 370574
rect 508266 334658 508502 334894
rect 508586 334658 508822 334894
rect 508266 334338 508502 334574
rect 508586 334338 508822 334574
rect 508266 298658 508502 298894
rect 508586 298658 508822 298894
rect 508266 298338 508502 298574
rect 508586 298338 508822 298574
rect 508266 262658 508502 262894
rect 508586 262658 508822 262894
rect 508266 262338 508502 262574
rect 508586 262338 508822 262574
rect 508266 226658 508502 226894
rect 508586 226658 508822 226894
rect 508266 226338 508502 226574
rect 508586 226338 508822 226574
rect 508266 190658 508502 190894
rect 508586 190658 508822 190894
rect 508266 190338 508502 190574
rect 508586 190338 508822 190574
rect 508266 154658 508502 154894
rect 508586 154658 508822 154894
rect 508266 154338 508502 154574
rect 508586 154338 508822 154574
rect 508266 118658 508502 118894
rect 508586 118658 508822 118894
rect 508266 118338 508502 118574
rect 508586 118338 508822 118574
rect 508266 82658 508502 82894
rect 508586 82658 508822 82894
rect 508266 82338 508502 82574
rect 508586 82338 508822 82574
rect 508266 46658 508502 46894
rect 508586 46658 508822 46894
rect 508266 46338 508502 46574
rect 508586 46338 508822 46574
rect 508266 10658 508502 10894
rect 508586 10658 508822 10894
rect 508266 10338 508502 10574
rect 508586 10338 508822 10574
rect 510826 705562 511062 705798
rect 511146 705562 511382 705798
rect 510826 705242 511062 705478
rect 511146 705242 511382 705478
rect 510826 669218 511062 669454
rect 511146 669218 511382 669454
rect 510826 668898 511062 669134
rect 511146 668898 511382 669134
rect 510826 633218 511062 633454
rect 511146 633218 511382 633454
rect 510826 632898 511062 633134
rect 511146 632898 511382 633134
rect 510826 597218 511062 597454
rect 511146 597218 511382 597454
rect 510826 596898 511062 597134
rect 511146 596898 511382 597134
rect 510826 561218 511062 561454
rect 511146 561218 511382 561454
rect 510826 560898 511062 561134
rect 511146 560898 511382 561134
rect 510826 525218 511062 525454
rect 511146 525218 511382 525454
rect 510826 524898 511062 525134
rect 511146 524898 511382 525134
rect 510826 489218 511062 489454
rect 511146 489218 511382 489454
rect 510826 488898 511062 489134
rect 511146 488898 511382 489134
rect 510826 453218 511062 453454
rect 511146 453218 511382 453454
rect 510826 452898 511062 453134
rect 511146 452898 511382 453134
rect 510826 417218 511062 417454
rect 511146 417218 511382 417454
rect 510826 416898 511062 417134
rect 511146 416898 511382 417134
rect 510826 381218 511062 381454
rect 511146 381218 511382 381454
rect 510826 380898 511062 381134
rect 511146 380898 511382 381134
rect 510826 345218 511062 345454
rect 511146 345218 511382 345454
rect 510826 344898 511062 345134
rect 511146 344898 511382 345134
rect 510826 309218 511062 309454
rect 511146 309218 511382 309454
rect 510826 308898 511062 309134
rect 511146 308898 511382 309134
rect 510826 273218 511062 273454
rect 511146 273218 511382 273454
rect 510826 272898 511062 273134
rect 511146 272898 511382 273134
rect 510826 237218 511062 237454
rect 511146 237218 511382 237454
rect 510826 236898 511062 237134
rect 511146 236898 511382 237134
rect 510826 201218 511062 201454
rect 511146 201218 511382 201454
rect 510826 200898 511062 201134
rect 511146 200898 511382 201134
rect 510826 165218 511062 165454
rect 511146 165218 511382 165454
rect 510826 164898 511062 165134
rect 511146 164898 511382 165134
rect 510826 129218 511062 129454
rect 511146 129218 511382 129454
rect 510826 128898 511062 129134
rect 511146 128898 511382 129134
rect 510826 93218 511062 93454
rect 511146 93218 511382 93454
rect 510826 92898 511062 93134
rect 511146 92898 511382 93134
rect 510826 57218 511062 57454
rect 511146 57218 511382 57454
rect 510826 56898 511062 57134
rect 511146 56898 511382 57134
rect 510826 21218 511062 21454
rect 511146 21218 511382 21454
rect 510826 20898 511062 21134
rect 511146 20898 511382 21134
rect 510826 -1542 511062 -1306
rect 511146 -1542 511382 -1306
rect 510826 -1862 511062 -1626
rect 511146 -1862 511382 -1626
rect 521986 711322 522222 711558
rect 522306 711322 522542 711558
rect 521986 711002 522222 711238
rect 522306 711002 522542 711238
rect 518266 709402 518502 709638
rect 518586 709402 518822 709638
rect 518266 709082 518502 709318
rect 518586 709082 518822 709318
rect 511986 698378 512222 698614
rect 512306 698378 512542 698614
rect 511986 698058 512222 698294
rect 512306 698058 512542 698294
rect 511986 662378 512222 662614
rect 512306 662378 512542 662614
rect 511986 662058 512222 662294
rect 512306 662058 512542 662294
rect 511986 626378 512222 626614
rect 512306 626378 512542 626614
rect 511986 626058 512222 626294
rect 512306 626058 512542 626294
rect 511986 590378 512222 590614
rect 512306 590378 512542 590614
rect 511986 590058 512222 590294
rect 512306 590058 512542 590294
rect 511986 554378 512222 554614
rect 512306 554378 512542 554614
rect 511986 554058 512222 554294
rect 512306 554058 512542 554294
rect 511986 518378 512222 518614
rect 512306 518378 512542 518614
rect 511986 518058 512222 518294
rect 512306 518058 512542 518294
rect 511986 482378 512222 482614
rect 512306 482378 512542 482614
rect 511986 482058 512222 482294
rect 512306 482058 512542 482294
rect 511986 446378 512222 446614
rect 512306 446378 512542 446614
rect 511986 446058 512222 446294
rect 512306 446058 512542 446294
rect 511986 410378 512222 410614
rect 512306 410378 512542 410614
rect 511986 410058 512222 410294
rect 512306 410058 512542 410294
rect 511986 374378 512222 374614
rect 512306 374378 512542 374614
rect 511986 374058 512222 374294
rect 512306 374058 512542 374294
rect 511986 338378 512222 338614
rect 512306 338378 512542 338614
rect 511986 338058 512222 338294
rect 512306 338058 512542 338294
rect 511986 302378 512222 302614
rect 512306 302378 512542 302614
rect 511986 302058 512222 302294
rect 512306 302058 512542 302294
rect 511986 266378 512222 266614
rect 512306 266378 512542 266614
rect 511986 266058 512222 266294
rect 512306 266058 512542 266294
rect 511986 230378 512222 230614
rect 512306 230378 512542 230614
rect 511986 230058 512222 230294
rect 512306 230058 512542 230294
rect 511986 194378 512222 194614
rect 512306 194378 512542 194614
rect 511986 194058 512222 194294
rect 512306 194058 512542 194294
rect 511986 158378 512222 158614
rect 512306 158378 512542 158614
rect 511986 158058 512222 158294
rect 512306 158058 512542 158294
rect 511986 122378 512222 122614
rect 512306 122378 512542 122614
rect 511986 122058 512222 122294
rect 512306 122058 512542 122294
rect 511986 86378 512222 86614
rect 512306 86378 512542 86614
rect 511986 86058 512222 86294
rect 512306 86058 512542 86294
rect 511986 50378 512222 50614
rect 512306 50378 512542 50614
rect 511986 50058 512222 50294
rect 512306 50058 512542 50294
rect 511986 14378 512222 14614
rect 512306 14378 512542 14614
rect 511986 14058 512222 14294
rect 512306 14058 512542 14294
rect 508266 -4422 508502 -4186
rect 508586 -4422 508822 -4186
rect 508266 -4742 508502 -4506
rect 508586 -4742 508822 -4506
rect 501986 -7302 502222 -7066
rect 502306 -7302 502542 -7066
rect 501986 -7622 502222 -7386
rect 502306 -7622 502542 -7386
rect 514546 707482 514782 707718
rect 514866 707482 515102 707718
rect 514546 707162 514782 707398
rect 514866 707162 515102 707398
rect 514546 672938 514782 673174
rect 514866 672938 515102 673174
rect 514546 672618 514782 672854
rect 514866 672618 515102 672854
rect 514546 636938 514782 637174
rect 514866 636938 515102 637174
rect 514546 636618 514782 636854
rect 514866 636618 515102 636854
rect 514546 600938 514782 601174
rect 514866 600938 515102 601174
rect 514546 600618 514782 600854
rect 514866 600618 515102 600854
rect 514546 564938 514782 565174
rect 514866 564938 515102 565174
rect 514546 564618 514782 564854
rect 514866 564618 515102 564854
rect 514546 528938 514782 529174
rect 514866 528938 515102 529174
rect 514546 528618 514782 528854
rect 514866 528618 515102 528854
rect 514546 492938 514782 493174
rect 514866 492938 515102 493174
rect 514546 492618 514782 492854
rect 514866 492618 515102 492854
rect 514546 456938 514782 457174
rect 514866 456938 515102 457174
rect 514546 456618 514782 456854
rect 514866 456618 515102 456854
rect 514546 420938 514782 421174
rect 514866 420938 515102 421174
rect 514546 420618 514782 420854
rect 514866 420618 515102 420854
rect 514546 384938 514782 385174
rect 514866 384938 515102 385174
rect 514546 384618 514782 384854
rect 514866 384618 515102 384854
rect 514546 348938 514782 349174
rect 514866 348938 515102 349174
rect 514546 348618 514782 348854
rect 514866 348618 515102 348854
rect 514546 312938 514782 313174
rect 514866 312938 515102 313174
rect 514546 312618 514782 312854
rect 514866 312618 515102 312854
rect 514546 276938 514782 277174
rect 514866 276938 515102 277174
rect 514546 276618 514782 276854
rect 514866 276618 515102 276854
rect 514546 240938 514782 241174
rect 514866 240938 515102 241174
rect 514546 240618 514782 240854
rect 514866 240618 515102 240854
rect 514546 204938 514782 205174
rect 514866 204938 515102 205174
rect 514546 204618 514782 204854
rect 514866 204618 515102 204854
rect 514546 168938 514782 169174
rect 514866 168938 515102 169174
rect 514546 168618 514782 168854
rect 514866 168618 515102 168854
rect 514546 132938 514782 133174
rect 514866 132938 515102 133174
rect 514546 132618 514782 132854
rect 514866 132618 515102 132854
rect 514546 96938 514782 97174
rect 514866 96938 515102 97174
rect 514546 96618 514782 96854
rect 514866 96618 515102 96854
rect 514546 60938 514782 61174
rect 514866 60938 515102 61174
rect 514546 60618 514782 60854
rect 514866 60618 515102 60854
rect 514546 24938 514782 25174
rect 514866 24938 515102 25174
rect 514546 24618 514782 24854
rect 514866 24618 515102 24854
rect 514546 -3462 514782 -3226
rect 514866 -3462 515102 -3226
rect 514546 -3782 514782 -3546
rect 514866 -3782 515102 -3546
rect 518266 676658 518502 676894
rect 518586 676658 518822 676894
rect 518266 676338 518502 676574
rect 518586 676338 518822 676574
rect 518266 640658 518502 640894
rect 518586 640658 518822 640894
rect 518266 640338 518502 640574
rect 518586 640338 518822 640574
rect 518266 604658 518502 604894
rect 518586 604658 518822 604894
rect 518266 604338 518502 604574
rect 518586 604338 518822 604574
rect 518266 568658 518502 568894
rect 518586 568658 518822 568894
rect 518266 568338 518502 568574
rect 518586 568338 518822 568574
rect 518266 532658 518502 532894
rect 518586 532658 518822 532894
rect 518266 532338 518502 532574
rect 518586 532338 518822 532574
rect 518266 496658 518502 496894
rect 518586 496658 518822 496894
rect 518266 496338 518502 496574
rect 518586 496338 518822 496574
rect 518266 460658 518502 460894
rect 518586 460658 518822 460894
rect 518266 460338 518502 460574
rect 518586 460338 518822 460574
rect 518266 424658 518502 424894
rect 518586 424658 518822 424894
rect 518266 424338 518502 424574
rect 518586 424338 518822 424574
rect 518266 388658 518502 388894
rect 518586 388658 518822 388894
rect 518266 388338 518502 388574
rect 518586 388338 518822 388574
rect 518266 352658 518502 352894
rect 518586 352658 518822 352894
rect 518266 352338 518502 352574
rect 518586 352338 518822 352574
rect 518266 316658 518502 316894
rect 518586 316658 518822 316894
rect 518266 316338 518502 316574
rect 518586 316338 518822 316574
rect 518266 280658 518502 280894
rect 518586 280658 518822 280894
rect 518266 280338 518502 280574
rect 518586 280338 518822 280574
rect 518266 244658 518502 244894
rect 518586 244658 518822 244894
rect 518266 244338 518502 244574
rect 518586 244338 518822 244574
rect 518266 208658 518502 208894
rect 518586 208658 518822 208894
rect 518266 208338 518502 208574
rect 518586 208338 518822 208574
rect 518266 172658 518502 172894
rect 518586 172658 518822 172894
rect 518266 172338 518502 172574
rect 518586 172338 518822 172574
rect 518266 136658 518502 136894
rect 518586 136658 518822 136894
rect 518266 136338 518502 136574
rect 518586 136338 518822 136574
rect 518266 100658 518502 100894
rect 518586 100658 518822 100894
rect 518266 100338 518502 100574
rect 518586 100338 518822 100574
rect 518266 64658 518502 64894
rect 518586 64658 518822 64894
rect 518266 64338 518502 64574
rect 518586 64338 518822 64574
rect 518266 28658 518502 28894
rect 518586 28658 518822 28894
rect 518266 28338 518502 28574
rect 518586 28338 518822 28574
rect 520826 704602 521062 704838
rect 521146 704602 521382 704838
rect 520826 704282 521062 704518
rect 521146 704282 521382 704518
rect 520826 687218 521062 687454
rect 521146 687218 521382 687454
rect 520826 686898 521062 687134
rect 521146 686898 521382 687134
rect 520826 651218 521062 651454
rect 521146 651218 521382 651454
rect 520826 650898 521062 651134
rect 521146 650898 521382 651134
rect 520826 615218 521062 615454
rect 521146 615218 521382 615454
rect 520826 614898 521062 615134
rect 521146 614898 521382 615134
rect 520826 579218 521062 579454
rect 521146 579218 521382 579454
rect 520826 578898 521062 579134
rect 521146 578898 521382 579134
rect 520826 543218 521062 543454
rect 521146 543218 521382 543454
rect 520826 542898 521062 543134
rect 521146 542898 521382 543134
rect 520826 507218 521062 507454
rect 521146 507218 521382 507454
rect 520826 506898 521062 507134
rect 521146 506898 521382 507134
rect 520826 471218 521062 471454
rect 521146 471218 521382 471454
rect 520826 470898 521062 471134
rect 521146 470898 521382 471134
rect 520826 435218 521062 435454
rect 521146 435218 521382 435454
rect 520826 434898 521062 435134
rect 521146 434898 521382 435134
rect 520826 399218 521062 399454
rect 521146 399218 521382 399454
rect 520826 398898 521062 399134
rect 521146 398898 521382 399134
rect 520826 363218 521062 363454
rect 521146 363218 521382 363454
rect 520826 362898 521062 363134
rect 521146 362898 521382 363134
rect 520826 327218 521062 327454
rect 521146 327218 521382 327454
rect 520826 326898 521062 327134
rect 521146 326898 521382 327134
rect 520826 291218 521062 291454
rect 521146 291218 521382 291454
rect 520826 290898 521062 291134
rect 521146 290898 521382 291134
rect 520826 255218 521062 255454
rect 521146 255218 521382 255454
rect 520826 254898 521062 255134
rect 521146 254898 521382 255134
rect 520826 219218 521062 219454
rect 521146 219218 521382 219454
rect 520826 218898 521062 219134
rect 521146 218898 521382 219134
rect 520826 183218 521062 183454
rect 521146 183218 521382 183454
rect 520826 182898 521062 183134
rect 521146 182898 521382 183134
rect 520826 147218 521062 147454
rect 521146 147218 521382 147454
rect 520826 146898 521062 147134
rect 521146 146898 521382 147134
rect 520826 111218 521062 111454
rect 521146 111218 521382 111454
rect 520826 110898 521062 111134
rect 521146 110898 521382 111134
rect 520826 75218 521062 75454
rect 521146 75218 521382 75454
rect 520826 74898 521062 75134
rect 521146 74898 521382 75134
rect 520826 39218 521062 39454
rect 521146 39218 521382 39454
rect 520826 38898 521062 39134
rect 521146 38898 521382 39134
rect 520826 3218 521062 3454
rect 521146 3218 521382 3454
rect 520826 2898 521062 3134
rect 521146 2898 521382 3134
rect 520826 -582 521062 -346
rect 521146 -582 521382 -346
rect 520826 -902 521062 -666
rect 521146 -902 521382 -666
rect 531986 710362 532222 710598
rect 532306 710362 532542 710598
rect 531986 710042 532222 710278
rect 532306 710042 532542 710278
rect 528266 708442 528502 708678
rect 528586 708442 528822 708678
rect 528266 708122 528502 708358
rect 528586 708122 528822 708358
rect 521986 680378 522222 680614
rect 522306 680378 522542 680614
rect 521986 680058 522222 680294
rect 522306 680058 522542 680294
rect 521986 644378 522222 644614
rect 522306 644378 522542 644614
rect 521986 644058 522222 644294
rect 522306 644058 522542 644294
rect 521986 608378 522222 608614
rect 522306 608378 522542 608614
rect 521986 608058 522222 608294
rect 522306 608058 522542 608294
rect 521986 572378 522222 572614
rect 522306 572378 522542 572614
rect 521986 572058 522222 572294
rect 522306 572058 522542 572294
rect 521986 536378 522222 536614
rect 522306 536378 522542 536614
rect 521986 536058 522222 536294
rect 522306 536058 522542 536294
rect 521986 500378 522222 500614
rect 522306 500378 522542 500614
rect 521986 500058 522222 500294
rect 522306 500058 522542 500294
rect 521986 464378 522222 464614
rect 522306 464378 522542 464614
rect 521986 464058 522222 464294
rect 522306 464058 522542 464294
rect 521986 428378 522222 428614
rect 522306 428378 522542 428614
rect 521986 428058 522222 428294
rect 522306 428058 522542 428294
rect 521986 392378 522222 392614
rect 522306 392378 522542 392614
rect 521986 392058 522222 392294
rect 522306 392058 522542 392294
rect 521986 356378 522222 356614
rect 522306 356378 522542 356614
rect 521986 356058 522222 356294
rect 522306 356058 522542 356294
rect 521986 320378 522222 320614
rect 522306 320378 522542 320614
rect 521986 320058 522222 320294
rect 522306 320058 522542 320294
rect 521986 284378 522222 284614
rect 522306 284378 522542 284614
rect 521986 284058 522222 284294
rect 522306 284058 522542 284294
rect 521986 248378 522222 248614
rect 522306 248378 522542 248614
rect 521986 248058 522222 248294
rect 522306 248058 522542 248294
rect 521986 212378 522222 212614
rect 522306 212378 522542 212614
rect 521986 212058 522222 212294
rect 522306 212058 522542 212294
rect 521986 176378 522222 176614
rect 522306 176378 522542 176614
rect 521986 176058 522222 176294
rect 522306 176058 522542 176294
rect 521986 140378 522222 140614
rect 522306 140378 522542 140614
rect 521986 140058 522222 140294
rect 522306 140058 522542 140294
rect 521986 104378 522222 104614
rect 522306 104378 522542 104614
rect 521986 104058 522222 104294
rect 522306 104058 522542 104294
rect 521986 68378 522222 68614
rect 522306 68378 522542 68614
rect 521986 68058 522222 68294
rect 522306 68058 522542 68294
rect 521986 32378 522222 32614
rect 522306 32378 522542 32614
rect 521986 32058 522222 32294
rect 522306 32058 522542 32294
rect 518266 -5382 518502 -5146
rect 518586 -5382 518822 -5146
rect 518266 -5702 518502 -5466
rect 518586 -5702 518822 -5466
rect 511986 -6342 512222 -6106
rect 512306 -6342 512542 -6106
rect 511986 -6662 512222 -6426
rect 512306 -6662 512542 -6426
rect 524546 706522 524782 706758
rect 524866 706522 525102 706758
rect 524546 706202 524782 706438
rect 524866 706202 525102 706438
rect 524546 690938 524782 691174
rect 524866 690938 525102 691174
rect 524546 690618 524782 690854
rect 524866 690618 525102 690854
rect 524546 654938 524782 655174
rect 524866 654938 525102 655174
rect 524546 654618 524782 654854
rect 524866 654618 525102 654854
rect 524546 618938 524782 619174
rect 524866 618938 525102 619174
rect 524546 618618 524782 618854
rect 524866 618618 525102 618854
rect 524546 582938 524782 583174
rect 524866 582938 525102 583174
rect 524546 582618 524782 582854
rect 524866 582618 525102 582854
rect 524546 546938 524782 547174
rect 524866 546938 525102 547174
rect 524546 546618 524782 546854
rect 524866 546618 525102 546854
rect 524546 510938 524782 511174
rect 524866 510938 525102 511174
rect 524546 510618 524782 510854
rect 524866 510618 525102 510854
rect 524546 474938 524782 475174
rect 524866 474938 525102 475174
rect 524546 474618 524782 474854
rect 524866 474618 525102 474854
rect 524546 438938 524782 439174
rect 524866 438938 525102 439174
rect 524546 438618 524782 438854
rect 524866 438618 525102 438854
rect 524546 402938 524782 403174
rect 524866 402938 525102 403174
rect 524546 402618 524782 402854
rect 524866 402618 525102 402854
rect 524546 366938 524782 367174
rect 524866 366938 525102 367174
rect 524546 366618 524782 366854
rect 524866 366618 525102 366854
rect 524546 330938 524782 331174
rect 524866 330938 525102 331174
rect 524546 330618 524782 330854
rect 524866 330618 525102 330854
rect 524546 294938 524782 295174
rect 524866 294938 525102 295174
rect 524546 294618 524782 294854
rect 524866 294618 525102 294854
rect 524546 258938 524782 259174
rect 524866 258938 525102 259174
rect 524546 258618 524782 258854
rect 524866 258618 525102 258854
rect 524546 222938 524782 223174
rect 524866 222938 525102 223174
rect 524546 222618 524782 222854
rect 524866 222618 525102 222854
rect 524546 186938 524782 187174
rect 524866 186938 525102 187174
rect 524546 186618 524782 186854
rect 524866 186618 525102 186854
rect 524546 150938 524782 151174
rect 524866 150938 525102 151174
rect 524546 150618 524782 150854
rect 524866 150618 525102 150854
rect 524546 114938 524782 115174
rect 524866 114938 525102 115174
rect 524546 114618 524782 114854
rect 524866 114618 525102 114854
rect 524546 78938 524782 79174
rect 524866 78938 525102 79174
rect 524546 78618 524782 78854
rect 524866 78618 525102 78854
rect 524546 42938 524782 43174
rect 524866 42938 525102 43174
rect 524546 42618 524782 42854
rect 524866 42618 525102 42854
rect 524546 6938 524782 7174
rect 524866 6938 525102 7174
rect 524546 6618 524782 6854
rect 524866 6618 525102 6854
rect 524546 -2502 524782 -2266
rect 524866 -2502 525102 -2266
rect 524546 -2822 524782 -2586
rect 524866 -2822 525102 -2586
rect 528266 694658 528502 694894
rect 528586 694658 528822 694894
rect 528266 694338 528502 694574
rect 528586 694338 528822 694574
rect 528266 658658 528502 658894
rect 528586 658658 528822 658894
rect 528266 658338 528502 658574
rect 528586 658338 528822 658574
rect 528266 622658 528502 622894
rect 528586 622658 528822 622894
rect 528266 622338 528502 622574
rect 528586 622338 528822 622574
rect 528266 586658 528502 586894
rect 528586 586658 528822 586894
rect 528266 586338 528502 586574
rect 528586 586338 528822 586574
rect 528266 550658 528502 550894
rect 528586 550658 528822 550894
rect 528266 550338 528502 550574
rect 528586 550338 528822 550574
rect 528266 514658 528502 514894
rect 528586 514658 528822 514894
rect 528266 514338 528502 514574
rect 528586 514338 528822 514574
rect 528266 478658 528502 478894
rect 528586 478658 528822 478894
rect 528266 478338 528502 478574
rect 528586 478338 528822 478574
rect 528266 442658 528502 442894
rect 528586 442658 528822 442894
rect 528266 442338 528502 442574
rect 528586 442338 528822 442574
rect 528266 406658 528502 406894
rect 528586 406658 528822 406894
rect 528266 406338 528502 406574
rect 528586 406338 528822 406574
rect 528266 370658 528502 370894
rect 528586 370658 528822 370894
rect 528266 370338 528502 370574
rect 528586 370338 528822 370574
rect 528266 334658 528502 334894
rect 528586 334658 528822 334894
rect 528266 334338 528502 334574
rect 528586 334338 528822 334574
rect 528266 298658 528502 298894
rect 528586 298658 528822 298894
rect 528266 298338 528502 298574
rect 528586 298338 528822 298574
rect 528266 262658 528502 262894
rect 528586 262658 528822 262894
rect 528266 262338 528502 262574
rect 528586 262338 528822 262574
rect 528266 226658 528502 226894
rect 528586 226658 528822 226894
rect 528266 226338 528502 226574
rect 528586 226338 528822 226574
rect 528266 190658 528502 190894
rect 528586 190658 528822 190894
rect 528266 190338 528502 190574
rect 528586 190338 528822 190574
rect 528266 154658 528502 154894
rect 528586 154658 528822 154894
rect 528266 154338 528502 154574
rect 528586 154338 528822 154574
rect 528266 118658 528502 118894
rect 528586 118658 528822 118894
rect 528266 118338 528502 118574
rect 528586 118338 528822 118574
rect 528266 82658 528502 82894
rect 528586 82658 528822 82894
rect 528266 82338 528502 82574
rect 528586 82338 528822 82574
rect 528266 46658 528502 46894
rect 528586 46658 528822 46894
rect 528266 46338 528502 46574
rect 528586 46338 528822 46574
rect 528266 10658 528502 10894
rect 528586 10658 528822 10894
rect 528266 10338 528502 10574
rect 528586 10338 528822 10574
rect 530826 705562 531062 705798
rect 531146 705562 531382 705798
rect 530826 705242 531062 705478
rect 531146 705242 531382 705478
rect 530826 669218 531062 669454
rect 531146 669218 531382 669454
rect 530826 668898 531062 669134
rect 531146 668898 531382 669134
rect 530826 633218 531062 633454
rect 531146 633218 531382 633454
rect 530826 632898 531062 633134
rect 531146 632898 531382 633134
rect 530826 597218 531062 597454
rect 531146 597218 531382 597454
rect 530826 596898 531062 597134
rect 531146 596898 531382 597134
rect 530826 561218 531062 561454
rect 531146 561218 531382 561454
rect 530826 560898 531062 561134
rect 531146 560898 531382 561134
rect 530826 525218 531062 525454
rect 531146 525218 531382 525454
rect 530826 524898 531062 525134
rect 531146 524898 531382 525134
rect 530826 489218 531062 489454
rect 531146 489218 531382 489454
rect 530826 488898 531062 489134
rect 531146 488898 531382 489134
rect 530826 453218 531062 453454
rect 531146 453218 531382 453454
rect 530826 452898 531062 453134
rect 531146 452898 531382 453134
rect 530826 417218 531062 417454
rect 531146 417218 531382 417454
rect 530826 416898 531062 417134
rect 531146 416898 531382 417134
rect 530826 381218 531062 381454
rect 531146 381218 531382 381454
rect 530826 380898 531062 381134
rect 531146 380898 531382 381134
rect 530826 345218 531062 345454
rect 531146 345218 531382 345454
rect 530826 344898 531062 345134
rect 531146 344898 531382 345134
rect 530826 309218 531062 309454
rect 531146 309218 531382 309454
rect 530826 308898 531062 309134
rect 531146 308898 531382 309134
rect 530826 273218 531062 273454
rect 531146 273218 531382 273454
rect 530826 272898 531062 273134
rect 531146 272898 531382 273134
rect 530826 237218 531062 237454
rect 531146 237218 531382 237454
rect 530826 236898 531062 237134
rect 531146 236898 531382 237134
rect 530826 201218 531062 201454
rect 531146 201218 531382 201454
rect 530826 200898 531062 201134
rect 531146 200898 531382 201134
rect 530826 165218 531062 165454
rect 531146 165218 531382 165454
rect 530826 164898 531062 165134
rect 531146 164898 531382 165134
rect 530826 129218 531062 129454
rect 531146 129218 531382 129454
rect 530826 128898 531062 129134
rect 531146 128898 531382 129134
rect 530826 93218 531062 93454
rect 531146 93218 531382 93454
rect 530826 92898 531062 93134
rect 531146 92898 531382 93134
rect 530826 57218 531062 57454
rect 531146 57218 531382 57454
rect 530826 56898 531062 57134
rect 531146 56898 531382 57134
rect 530826 21218 531062 21454
rect 531146 21218 531382 21454
rect 530826 20898 531062 21134
rect 531146 20898 531382 21134
rect 530826 -1542 531062 -1306
rect 531146 -1542 531382 -1306
rect 530826 -1862 531062 -1626
rect 531146 -1862 531382 -1626
rect 541986 711322 542222 711558
rect 542306 711322 542542 711558
rect 541986 711002 542222 711238
rect 542306 711002 542542 711238
rect 538266 709402 538502 709638
rect 538586 709402 538822 709638
rect 538266 709082 538502 709318
rect 538586 709082 538822 709318
rect 531986 698378 532222 698614
rect 532306 698378 532542 698614
rect 531986 698058 532222 698294
rect 532306 698058 532542 698294
rect 531986 662378 532222 662614
rect 532306 662378 532542 662614
rect 531986 662058 532222 662294
rect 532306 662058 532542 662294
rect 531986 626378 532222 626614
rect 532306 626378 532542 626614
rect 531986 626058 532222 626294
rect 532306 626058 532542 626294
rect 531986 590378 532222 590614
rect 532306 590378 532542 590614
rect 531986 590058 532222 590294
rect 532306 590058 532542 590294
rect 531986 554378 532222 554614
rect 532306 554378 532542 554614
rect 531986 554058 532222 554294
rect 532306 554058 532542 554294
rect 531986 518378 532222 518614
rect 532306 518378 532542 518614
rect 531986 518058 532222 518294
rect 532306 518058 532542 518294
rect 531986 482378 532222 482614
rect 532306 482378 532542 482614
rect 531986 482058 532222 482294
rect 532306 482058 532542 482294
rect 531986 446378 532222 446614
rect 532306 446378 532542 446614
rect 531986 446058 532222 446294
rect 532306 446058 532542 446294
rect 531986 410378 532222 410614
rect 532306 410378 532542 410614
rect 531986 410058 532222 410294
rect 532306 410058 532542 410294
rect 531986 374378 532222 374614
rect 532306 374378 532542 374614
rect 531986 374058 532222 374294
rect 532306 374058 532542 374294
rect 531986 338378 532222 338614
rect 532306 338378 532542 338614
rect 531986 338058 532222 338294
rect 532306 338058 532542 338294
rect 531986 302378 532222 302614
rect 532306 302378 532542 302614
rect 531986 302058 532222 302294
rect 532306 302058 532542 302294
rect 531986 266378 532222 266614
rect 532306 266378 532542 266614
rect 531986 266058 532222 266294
rect 532306 266058 532542 266294
rect 531986 230378 532222 230614
rect 532306 230378 532542 230614
rect 531986 230058 532222 230294
rect 532306 230058 532542 230294
rect 531986 194378 532222 194614
rect 532306 194378 532542 194614
rect 531986 194058 532222 194294
rect 532306 194058 532542 194294
rect 531986 158378 532222 158614
rect 532306 158378 532542 158614
rect 531986 158058 532222 158294
rect 532306 158058 532542 158294
rect 531986 122378 532222 122614
rect 532306 122378 532542 122614
rect 531986 122058 532222 122294
rect 532306 122058 532542 122294
rect 531986 86378 532222 86614
rect 532306 86378 532542 86614
rect 531986 86058 532222 86294
rect 532306 86058 532542 86294
rect 531986 50378 532222 50614
rect 532306 50378 532542 50614
rect 531986 50058 532222 50294
rect 532306 50058 532542 50294
rect 531986 14378 532222 14614
rect 532306 14378 532542 14614
rect 531986 14058 532222 14294
rect 532306 14058 532542 14294
rect 528266 -4422 528502 -4186
rect 528586 -4422 528822 -4186
rect 528266 -4742 528502 -4506
rect 528586 -4742 528822 -4506
rect 521986 -7302 522222 -7066
rect 522306 -7302 522542 -7066
rect 521986 -7622 522222 -7386
rect 522306 -7622 522542 -7386
rect 534546 707482 534782 707718
rect 534866 707482 535102 707718
rect 534546 707162 534782 707398
rect 534866 707162 535102 707398
rect 534546 672938 534782 673174
rect 534866 672938 535102 673174
rect 534546 672618 534782 672854
rect 534866 672618 535102 672854
rect 534546 636938 534782 637174
rect 534866 636938 535102 637174
rect 534546 636618 534782 636854
rect 534866 636618 535102 636854
rect 534546 600938 534782 601174
rect 534866 600938 535102 601174
rect 534546 600618 534782 600854
rect 534866 600618 535102 600854
rect 534546 564938 534782 565174
rect 534866 564938 535102 565174
rect 534546 564618 534782 564854
rect 534866 564618 535102 564854
rect 534546 528938 534782 529174
rect 534866 528938 535102 529174
rect 534546 528618 534782 528854
rect 534866 528618 535102 528854
rect 534546 492938 534782 493174
rect 534866 492938 535102 493174
rect 534546 492618 534782 492854
rect 534866 492618 535102 492854
rect 534546 456938 534782 457174
rect 534866 456938 535102 457174
rect 534546 456618 534782 456854
rect 534866 456618 535102 456854
rect 534546 420938 534782 421174
rect 534866 420938 535102 421174
rect 534546 420618 534782 420854
rect 534866 420618 535102 420854
rect 534546 384938 534782 385174
rect 534866 384938 535102 385174
rect 534546 384618 534782 384854
rect 534866 384618 535102 384854
rect 534546 348938 534782 349174
rect 534866 348938 535102 349174
rect 534546 348618 534782 348854
rect 534866 348618 535102 348854
rect 534546 312938 534782 313174
rect 534866 312938 535102 313174
rect 534546 312618 534782 312854
rect 534866 312618 535102 312854
rect 534546 276938 534782 277174
rect 534866 276938 535102 277174
rect 534546 276618 534782 276854
rect 534866 276618 535102 276854
rect 534546 240938 534782 241174
rect 534866 240938 535102 241174
rect 534546 240618 534782 240854
rect 534866 240618 535102 240854
rect 534546 204938 534782 205174
rect 534866 204938 535102 205174
rect 534546 204618 534782 204854
rect 534866 204618 535102 204854
rect 534546 168938 534782 169174
rect 534866 168938 535102 169174
rect 534546 168618 534782 168854
rect 534866 168618 535102 168854
rect 534546 132938 534782 133174
rect 534866 132938 535102 133174
rect 534546 132618 534782 132854
rect 534866 132618 535102 132854
rect 534546 96938 534782 97174
rect 534866 96938 535102 97174
rect 534546 96618 534782 96854
rect 534866 96618 535102 96854
rect 534546 60938 534782 61174
rect 534866 60938 535102 61174
rect 534546 60618 534782 60854
rect 534866 60618 535102 60854
rect 534546 24938 534782 25174
rect 534866 24938 535102 25174
rect 534546 24618 534782 24854
rect 534866 24618 535102 24854
rect 534546 -3462 534782 -3226
rect 534866 -3462 535102 -3226
rect 534546 -3782 534782 -3546
rect 534866 -3782 535102 -3546
rect 538266 676658 538502 676894
rect 538586 676658 538822 676894
rect 538266 676338 538502 676574
rect 538586 676338 538822 676574
rect 538266 640658 538502 640894
rect 538586 640658 538822 640894
rect 538266 640338 538502 640574
rect 538586 640338 538822 640574
rect 538266 604658 538502 604894
rect 538586 604658 538822 604894
rect 538266 604338 538502 604574
rect 538586 604338 538822 604574
rect 538266 568658 538502 568894
rect 538586 568658 538822 568894
rect 538266 568338 538502 568574
rect 538586 568338 538822 568574
rect 538266 532658 538502 532894
rect 538586 532658 538822 532894
rect 538266 532338 538502 532574
rect 538586 532338 538822 532574
rect 538266 496658 538502 496894
rect 538586 496658 538822 496894
rect 538266 496338 538502 496574
rect 538586 496338 538822 496574
rect 538266 460658 538502 460894
rect 538586 460658 538822 460894
rect 538266 460338 538502 460574
rect 538586 460338 538822 460574
rect 538266 424658 538502 424894
rect 538586 424658 538822 424894
rect 538266 424338 538502 424574
rect 538586 424338 538822 424574
rect 538266 388658 538502 388894
rect 538586 388658 538822 388894
rect 538266 388338 538502 388574
rect 538586 388338 538822 388574
rect 538266 352658 538502 352894
rect 538586 352658 538822 352894
rect 538266 352338 538502 352574
rect 538586 352338 538822 352574
rect 538266 316658 538502 316894
rect 538586 316658 538822 316894
rect 538266 316338 538502 316574
rect 538586 316338 538822 316574
rect 538266 280658 538502 280894
rect 538586 280658 538822 280894
rect 538266 280338 538502 280574
rect 538586 280338 538822 280574
rect 538266 244658 538502 244894
rect 538586 244658 538822 244894
rect 538266 244338 538502 244574
rect 538586 244338 538822 244574
rect 538266 208658 538502 208894
rect 538586 208658 538822 208894
rect 538266 208338 538502 208574
rect 538586 208338 538822 208574
rect 538266 172658 538502 172894
rect 538586 172658 538822 172894
rect 538266 172338 538502 172574
rect 538586 172338 538822 172574
rect 538266 136658 538502 136894
rect 538586 136658 538822 136894
rect 538266 136338 538502 136574
rect 538586 136338 538822 136574
rect 538266 100658 538502 100894
rect 538586 100658 538822 100894
rect 538266 100338 538502 100574
rect 538586 100338 538822 100574
rect 538266 64658 538502 64894
rect 538586 64658 538822 64894
rect 538266 64338 538502 64574
rect 538586 64338 538822 64574
rect 538266 28658 538502 28894
rect 538586 28658 538822 28894
rect 538266 28338 538502 28574
rect 538586 28338 538822 28574
rect 540826 704602 541062 704838
rect 541146 704602 541382 704838
rect 540826 704282 541062 704518
rect 541146 704282 541382 704518
rect 540826 687218 541062 687454
rect 541146 687218 541382 687454
rect 540826 686898 541062 687134
rect 541146 686898 541382 687134
rect 540826 651218 541062 651454
rect 541146 651218 541382 651454
rect 540826 650898 541062 651134
rect 541146 650898 541382 651134
rect 540826 615218 541062 615454
rect 541146 615218 541382 615454
rect 540826 614898 541062 615134
rect 541146 614898 541382 615134
rect 540826 579218 541062 579454
rect 541146 579218 541382 579454
rect 540826 578898 541062 579134
rect 541146 578898 541382 579134
rect 540826 543218 541062 543454
rect 541146 543218 541382 543454
rect 540826 542898 541062 543134
rect 541146 542898 541382 543134
rect 540826 507218 541062 507454
rect 541146 507218 541382 507454
rect 540826 506898 541062 507134
rect 541146 506898 541382 507134
rect 540826 471218 541062 471454
rect 541146 471218 541382 471454
rect 540826 470898 541062 471134
rect 541146 470898 541382 471134
rect 540826 435218 541062 435454
rect 541146 435218 541382 435454
rect 540826 434898 541062 435134
rect 541146 434898 541382 435134
rect 540826 399218 541062 399454
rect 541146 399218 541382 399454
rect 540826 398898 541062 399134
rect 541146 398898 541382 399134
rect 540826 363218 541062 363454
rect 541146 363218 541382 363454
rect 540826 362898 541062 363134
rect 541146 362898 541382 363134
rect 540826 327218 541062 327454
rect 541146 327218 541382 327454
rect 540826 326898 541062 327134
rect 541146 326898 541382 327134
rect 540826 291218 541062 291454
rect 541146 291218 541382 291454
rect 540826 290898 541062 291134
rect 541146 290898 541382 291134
rect 540826 255218 541062 255454
rect 541146 255218 541382 255454
rect 540826 254898 541062 255134
rect 541146 254898 541382 255134
rect 540826 219218 541062 219454
rect 541146 219218 541382 219454
rect 540826 218898 541062 219134
rect 541146 218898 541382 219134
rect 540826 183218 541062 183454
rect 541146 183218 541382 183454
rect 540826 182898 541062 183134
rect 541146 182898 541382 183134
rect 540826 147218 541062 147454
rect 541146 147218 541382 147454
rect 540826 146898 541062 147134
rect 541146 146898 541382 147134
rect 540826 111218 541062 111454
rect 541146 111218 541382 111454
rect 540826 110898 541062 111134
rect 541146 110898 541382 111134
rect 540826 75218 541062 75454
rect 541146 75218 541382 75454
rect 540826 74898 541062 75134
rect 541146 74898 541382 75134
rect 540826 39218 541062 39454
rect 541146 39218 541382 39454
rect 540826 38898 541062 39134
rect 541146 38898 541382 39134
rect 540826 3218 541062 3454
rect 541146 3218 541382 3454
rect 540826 2898 541062 3134
rect 541146 2898 541382 3134
rect 540826 -582 541062 -346
rect 541146 -582 541382 -346
rect 540826 -902 541062 -666
rect 541146 -902 541382 -666
rect 551986 710362 552222 710598
rect 552306 710362 552542 710598
rect 551986 710042 552222 710278
rect 552306 710042 552542 710278
rect 548266 708442 548502 708678
rect 548586 708442 548822 708678
rect 548266 708122 548502 708358
rect 548586 708122 548822 708358
rect 541986 680378 542222 680614
rect 542306 680378 542542 680614
rect 541986 680058 542222 680294
rect 542306 680058 542542 680294
rect 541986 644378 542222 644614
rect 542306 644378 542542 644614
rect 541986 644058 542222 644294
rect 542306 644058 542542 644294
rect 541986 608378 542222 608614
rect 542306 608378 542542 608614
rect 541986 608058 542222 608294
rect 542306 608058 542542 608294
rect 541986 572378 542222 572614
rect 542306 572378 542542 572614
rect 541986 572058 542222 572294
rect 542306 572058 542542 572294
rect 541986 536378 542222 536614
rect 542306 536378 542542 536614
rect 541986 536058 542222 536294
rect 542306 536058 542542 536294
rect 541986 500378 542222 500614
rect 542306 500378 542542 500614
rect 541986 500058 542222 500294
rect 542306 500058 542542 500294
rect 541986 464378 542222 464614
rect 542306 464378 542542 464614
rect 541986 464058 542222 464294
rect 542306 464058 542542 464294
rect 541986 428378 542222 428614
rect 542306 428378 542542 428614
rect 541986 428058 542222 428294
rect 542306 428058 542542 428294
rect 541986 392378 542222 392614
rect 542306 392378 542542 392614
rect 541986 392058 542222 392294
rect 542306 392058 542542 392294
rect 541986 356378 542222 356614
rect 542306 356378 542542 356614
rect 541986 356058 542222 356294
rect 542306 356058 542542 356294
rect 541986 320378 542222 320614
rect 542306 320378 542542 320614
rect 541986 320058 542222 320294
rect 542306 320058 542542 320294
rect 541986 284378 542222 284614
rect 542306 284378 542542 284614
rect 541986 284058 542222 284294
rect 542306 284058 542542 284294
rect 541986 248378 542222 248614
rect 542306 248378 542542 248614
rect 541986 248058 542222 248294
rect 542306 248058 542542 248294
rect 541986 212378 542222 212614
rect 542306 212378 542542 212614
rect 541986 212058 542222 212294
rect 542306 212058 542542 212294
rect 541986 176378 542222 176614
rect 542306 176378 542542 176614
rect 541986 176058 542222 176294
rect 542306 176058 542542 176294
rect 541986 140378 542222 140614
rect 542306 140378 542542 140614
rect 541986 140058 542222 140294
rect 542306 140058 542542 140294
rect 541986 104378 542222 104614
rect 542306 104378 542542 104614
rect 541986 104058 542222 104294
rect 542306 104058 542542 104294
rect 541986 68378 542222 68614
rect 542306 68378 542542 68614
rect 541986 68058 542222 68294
rect 542306 68058 542542 68294
rect 541986 32378 542222 32614
rect 542306 32378 542542 32614
rect 541986 32058 542222 32294
rect 542306 32058 542542 32294
rect 538266 -5382 538502 -5146
rect 538586 -5382 538822 -5146
rect 538266 -5702 538502 -5466
rect 538586 -5702 538822 -5466
rect 531986 -6342 532222 -6106
rect 532306 -6342 532542 -6106
rect 531986 -6662 532222 -6426
rect 532306 -6662 532542 -6426
rect 544546 706522 544782 706758
rect 544866 706522 545102 706758
rect 544546 706202 544782 706438
rect 544866 706202 545102 706438
rect 544546 690938 544782 691174
rect 544866 690938 545102 691174
rect 544546 690618 544782 690854
rect 544866 690618 545102 690854
rect 544546 654938 544782 655174
rect 544866 654938 545102 655174
rect 544546 654618 544782 654854
rect 544866 654618 545102 654854
rect 544546 618938 544782 619174
rect 544866 618938 545102 619174
rect 544546 618618 544782 618854
rect 544866 618618 545102 618854
rect 544546 582938 544782 583174
rect 544866 582938 545102 583174
rect 544546 582618 544782 582854
rect 544866 582618 545102 582854
rect 544546 546938 544782 547174
rect 544866 546938 545102 547174
rect 544546 546618 544782 546854
rect 544866 546618 545102 546854
rect 544546 510938 544782 511174
rect 544866 510938 545102 511174
rect 544546 510618 544782 510854
rect 544866 510618 545102 510854
rect 544546 474938 544782 475174
rect 544866 474938 545102 475174
rect 544546 474618 544782 474854
rect 544866 474618 545102 474854
rect 544546 438938 544782 439174
rect 544866 438938 545102 439174
rect 544546 438618 544782 438854
rect 544866 438618 545102 438854
rect 544546 402938 544782 403174
rect 544866 402938 545102 403174
rect 544546 402618 544782 402854
rect 544866 402618 545102 402854
rect 544546 366938 544782 367174
rect 544866 366938 545102 367174
rect 544546 366618 544782 366854
rect 544866 366618 545102 366854
rect 544546 330938 544782 331174
rect 544866 330938 545102 331174
rect 544546 330618 544782 330854
rect 544866 330618 545102 330854
rect 544546 294938 544782 295174
rect 544866 294938 545102 295174
rect 544546 294618 544782 294854
rect 544866 294618 545102 294854
rect 544546 258938 544782 259174
rect 544866 258938 545102 259174
rect 544546 258618 544782 258854
rect 544866 258618 545102 258854
rect 544546 222938 544782 223174
rect 544866 222938 545102 223174
rect 544546 222618 544782 222854
rect 544866 222618 545102 222854
rect 544546 186938 544782 187174
rect 544866 186938 545102 187174
rect 544546 186618 544782 186854
rect 544866 186618 545102 186854
rect 544546 150938 544782 151174
rect 544866 150938 545102 151174
rect 544546 150618 544782 150854
rect 544866 150618 545102 150854
rect 544546 114938 544782 115174
rect 544866 114938 545102 115174
rect 544546 114618 544782 114854
rect 544866 114618 545102 114854
rect 544546 78938 544782 79174
rect 544866 78938 545102 79174
rect 544546 78618 544782 78854
rect 544866 78618 545102 78854
rect 544546 42938 544782 43174
rect 544866 42938 545102 43174
rect 544546 42618 544782 42854
rect 544866 42618 545102 42854
rect 544546 6938 544782 7174
rect 544866 6938 545102 7174
rect 544546 6618 544782 6854
rect 544866 6618 545102 6854
rect 544546 -2502 544782 -2266
rect 544866 -2502 545102 -2266
rect 544546 -2822 544782 -2586
rect 544866 -2822 545102 -2586
rect 548266 694658 548502 694894
rect 548586 694658 548822 694894
rect 548266 694338 548502 694574
rect 548586 694338 548822 694574
rect 548266 658658 548502 658894
rect 548586 658658 548822 658894
rect 548266 658338 548502 658574
rect 548586 658338 548822 658574
rect 548266 622658 548502 622894
rect 548586 622658 548822 622894
rect 548266 622338 548502 622574
rect 548586 622338 548822 622574
rect 548266 586658 548502 586894
rect 548586 586658 548822 586894
rect 548266 586338 548502 586574
rect 548586 586338 548822 586574
rect 548266 550658 548502 550894
rect 548586 550658 548822 550894
rect 548266 550338 548502 550574
rect 548586 550338 548822 550574
rect 548266 514658 548502 514894
rect 548586 514658 548822 514894
rect 548266 514338 548502 514574
rect 548586 514338 548822 514574
rect 548266 478658 548502 478894
rect 548586 478658 548822 478894
rect 548266 478338 548502 478574
rect 548586 478338 548822 478574
rect 548266 442658 548502 442894
rect 548586 442658 548822 442894
rect 548266 442338 548502 442574
rect 548586 442338 548822 442574
rect 548266 406658 548502 406894
rect 548586 406658 548822 406894
rect 548266 406338 548502 406574
rect 548586 406338 548822 406574
rect 548266 370658 548502 370894
rect 548586 370658 548822 370894
rect 548266 370338 548502 370574
rect 548586 370338 548822 370574
rect 548266 334658 548502 334894
rect 548586 334658 548822 334894
rect 548266 334338 548502 334574
rect 548586 334338 548822 334574
rect 548266 298658 548502 298894
rect 548586 298658 548822 298894
rect 548266 298338 548502 298574
rect 548586 298338 548822 298574
rect 548266 262658 548502 262894
rect 548586 262658 548822 262894
rect 548266 262338 548502 262574
rect 548586 262338 548822 262574
rect 548266 226658 548502 226894
rect 548586 226658 548822 226894
rect 548266 226338 548502 226574
rect 548586 226338 548822 226574
rect 548266 190658 548502 190894
rect 548586 190658 548822 190894
rect 548266 190338 548502 190574
rect 548586 190338 548822 190574
rect 548266 154658 548502 154894
rect 548586 154658 548822 154894
rect 548266 154338 548502 154574
rect 548586 154338 548822 154574
rect 548266 118658 548502 118894
rect 548586 118658 548822 118894
rect 548266 118338 548502 118574
rect 548586 118338 548822 118574
rect 548266 82658 548502 82894
rect 548586 82658 548822 82894
rect 548266 82338 548502 82574
rect 548586 82338 548822 82574
rect 548266 46658 548502 46894
rect 548586 46658 548822 46894
rect 548266 46338 548502 46574
rect 548586 46338 548822 46574
rect 548266 10658 548502 10894
rect 548586 10658 548822 10894
rect 548266 10338 548502 10574
rect 548586 10338 548822 10574
rect 550826 705562 551062 705798
rect 551146 705562 551382 705798
rect 550826 705242 551062 705478
rect 551146 705242 551382 705478
rect 550826 669218 551062 669454
rect 551146 669218 551382 669454
rect 550826 668898 551062 669134
rect 551146 668898 551382 669134
rect 550826 633218 551062 633454
rect 551146 633218 551382 633454
rect 550826 632898 551062 633134
rect 551146 632898 551382 633134
rect 550826 597218 551062 597454
rect 551146 597218 551382 597454
rect 550826 596898 551062 597134
rect 551146 596898 551382 597134
rect 550826 561218 551062 561454
rect 551146 561218 551382 561454
rect 550826 560898 551062 561134
rect 551146 560898 551382 561134
rect 550826 525218 551062 525454
rect 551146 525218 551382 525454
rect 550826 524898 551062 525134
rect 551146 524898 551382 525134
rect 550826 489218 551062 489454
rect 551146 489218 551382 489454
rect 550826 488898 551062 489134
rect 551146 488898 551382 489134
rect 550826 453218 551062 453454
rect 551146 453218 551382 453454
rect 550826 452898 551062 453134
rect 551146 452898 551382 453134
rect 550826 417218 551062 417454
rect 551146 417218 551382 417454
rect 550826 416898 551062 417134
rect 551146 416898 551382 417134
rect 550826 381218 551062 381454
rect 551146 381218 551382 381454
rect 550826 380898 551062 381134
rect 551146 380898 551382 381134
rect 550826 345218 551062 345454
rect 551146 345218 551382 345454
rect 550826 344898 551062 345134
rect 551146 344898 551382 345134
rect 550826 309218 551062 309454
rect 551146 309218 551382 309454
rect 550826 308898 551062 309134
rect 551146 308898 551382 309134
rect 550826 273218 551062 273454
rect 551146 273218 551382 273454
rect 550826 272898 551062 273134
rect 551146 272898 551382 273134
rect 550826 237218 551062 237454
rect 551146 237218 551382 237454
rect 550826 236898 551062 237134
rect 551146 236898 551382 237134
rect 550826 201218 551062 201454
rect 551146 201218 551382 201454
rect 550826 200898 551062 201134
rect 551146 200898 551382 201134
rect 550826 165218 551062 165454
rect 551146 165218 551382 165454
rect 550826 164898 551062 165134
rect 551146 164898 551382 165134
rect 550826 129218 551062 129454
rect 551146 129218 551382 129454
rect 550826 128898 551062 129134
rect 551146 128898 551382 129134
rect 550826 93218 551062 93454
rect 551146 93218 551382 93454
rect 550826 92898 551062 93134
rect 551146 92898 551382 93134
rect 550826 57218 551062 57454
rect 551146 57218 551382 57454
rect 550826 56898 551062 57134
rect 551146 56898 551382 57134
rect 550826 21218 551062 21454
rect 551146 21218 551382 21454
rect 550826 20898 551062 21134
rect 551146 20898 551382 21134
rect 550826 -1542 551062 -1306
rect 551146 -1542 551382 -1306
rect 550826 -1862 551062 -1626
rect 551146 -1862 551382 -1626
rect 561986 711322 562222 711558
rect 562306 711322 562542 711558
rect 561986 711002 562222 711238
rect 562306 711002 562542 711238
rect 558266 709402 558502 709638
rect 558586 709402 558822 709638
rect 558266 709082 558502 709318
rect 558586 709082 558822 709318
rect 551986 698378 552222 698614
rect 552306 698378 552542 698614
rect 551986 698058 552222 698294
rect 552306 698058 552542 698294
rect 551986 662378 552222 662614
rect 552306 662378 552542 662614
rect 551986 662058 552222 662294
rect 552306 662058 552542 662294
rect 551986 626378 552222 626614
rect 552306 626378 552542 626614
rect 551986 626058 552222 626294
rect 552306 626058 552542 626294
rect 551986 590378 552222 590614
rect 552306 590378 552542 590614
rect 551986 590058 552222 590294
rect 552306 590058 552542 590294
rect 551986 554378 552222 554614
rect 552306 554378 552542 554614
rect 551986 554058 552222 554294
rect 552306 554058 552542 554294
rect 551986 518378 552222 518614
rect 552306 518378 552542 518614
rect 551986 518058 552222 518294
rect 552306 518058 552542 518294
rect 551986 482378 552222 482614
rect 552306 482378 552542 482614
rect 551986 482058 552222 482294
rect 552306 482058 552542 482294
rect 551986 446378 552222 446614
rect 552306 446378 552542 446614
rect 551986 446058 552222 446294
rect 552306 446058 552542 446294
rect 551986 410378 552222 410614
rect 552306 410378 552542 410614
rect 551986 410058 552222 410294
rect 552306 410058 552542 410294
rect 551986 374378 552222 374614
rect 552306 374378 552542 374614
rect 551986 374058 552222 374294
rect 552306 374058 552542 374294
rect 551986 338378 552222 338614
rect 552306 338378 552542 338614
rect 551986 338058 552222 338294
rect 552306 338058 552542 338294
rect 551986 302378 552222 302614
rect 552306 302378 552542 302614
rect 551986 302058 552222 302294
rect 552306 302058 552542 302294
rect 551986 266378 552222 266614
rect 552306 266378 552542 266614
rect 551986 266058 552222 266294
rect 552306 266058 552542 266294
rect 551986 230378 552222 230614
rect 552306 230378 552542 230614
rect 551986 230058 552222 230294
rect 552306 230058 552542 230294
rect 551986 194378 552222 194614
rect 552306 194378 552542 194614
rect 551986 194058 552222 194294
rect 552306 194058 552542 194294
rect 551986 158378 552222 158614
rect 552306 158378 552542 158614
rect 551986 158058 552222 158294
rect 552306 158058 552542 158294
rect 551986 122378 552222 122614
rect 552306 122378 552542 122614
rect 551986 122058 552222 122294
rect 552306 122058 552542 122294
rect 551986 86378 552222 86614
rect 552306 86378 552542 86614
rect 551986 86058 552222 86294
rect 552306 86058 552542 86294
rect 551986 50378 552222 50614
rect 552306 50378 552542 50614
rect 551986 50058 552222 50294
rect 552306 50058 552542 50294
rect 551986 14378 552222 14614
rect 552306 14378 552542 14614
rect 551986 14058 552222 14294
rect 552306 14058 552542 14294
rect 548266 -4422 548502 -4186
rect 548586 -4422 548822 -4186
rect 548266 -4742 548502 -4506
rect 548586 -4742 548822 -4506
rect 541986 -7302 542222 -7066
rect 542306 -7302 542542 -7066
rect 541986 -7622 542222 -7386
rect 542306 -7622 542542 -7386
rect 554546 707482 554782 707718
rect 554866 707482 555102 707718
rect 554546 707162 554782 707398
rect 554866 707162 555102 707398
rect 554546 672938 554782 673174
rect 554866 672938 555102 673174
rect 554546 672618 554782 672854
rect 554866 672618 555102 672854
rect 554546 636938 554782 637174
rect 554866 636938 555102 637174
rect 554546 636618 554782 636854
rect 554866 636618 555102 636854
rect 554546 600938 554782 601174
rect 554866 600938 555102 601174
rect 554546 600618 554782 600854
rect 554866 600618 555102 600854
rect 554546 564938 554782 565174
rect 554866 564938 555102 565174
rect 554546 564618 554782 564854
rect 554866 564618 555102 564854
rect 554546 528938 554782 529174
rect 554866 528938 555102 529174
rect 554546 528618 554782 528854
rect 554866 528618 555102 528854
rect 554546 492938 554782 493174
rect 554866 492938 555102 493174
rect 554546 492618 554782 492854
rect 554866 492618 555102 492854
rect 554546 456938 554782 457174
rect 554866 456938 555102 457174
rect 554546 456618 554782 456854
rect 554866 456618 555102 456854
rect 554546 420938 554782 421174
rect 554866 420938 555102 421174
rect 554546 420618 554782 420854
rect 554866 420618 555102 420854
rect 554546 384938 554782 385174
rect 554866 384938 555102 385174
rect 554546 384618 554782 384854
rect 554866 384618 555102 384854
rect 554546 348938 554782 349174
rect 554866 348938 555102 349174
rect 554546 348618 554782 348854
rect 554866 348618 555102 348854
rect 554546 312938 554782 313174
rect 554866 312938 555102 313174
rect 554546 312618 554782 312854
rect 554866 312618 555102 312854
rect 554546 276938 554782 277174
rect 554866 276938 555102 277174
rect 554546 276618 554782 276854
rect 554866 276618 555102 276854
rect 554546 240938 554782 241174
rect 554866 240938 555102 241174
rect 554546 240618 554782 240854
rect 554866 240618 555102 240854
rect 554546 204938 554782 205174
rect 554866 204938 555102 205174
rect 554546 204618 554782 204854
rect 554866 204618 555102 204854
rect 554546 168938 554782 169174
rect 554866 168938 555102 169174
rect 554546 168618 554782 168854
rect 554866 168618 555102 168854
rect 554546 132938 554782 133174
rect 554866 132938 555102 133174
rect 554546 132618 554782 132854
rect 554866 132618 555102 132854
rect 554546 96938 554782 97174
rect 554866 96938 555102 97174
rect 554546 96618 554782 96854
rect 554866 96618 555102 96854
rect 554546 60938 554782 61174
rect 554866 60938 555102 61174
rect 554546 60618 554782 60854
rect 554866 60618 555102 60854
rect 554546 24938 554782 25174
rect 554866 24938 555102 25174
rect 554546 24618 554782 24854
rect 554866 24618 555102 24854
rect 554546 -3462 554782 -3226
rect 554866 -3462 555102 -3226
rect 554546 -3782 554782 -3546
rect 554866 -3782 555102 -3546
rect 558266 676658 558502 676894
rect 558586 676658 558822 676894
rect 558266 676338 558502 676574
rect 558586 676338 558822 676574
rect 558266 640658 558502 640894
rect 558586 640658 558822 640894
rect 558266 640338 558502 640574
rect 558586 640338 558822 640574
rect 558266 604658 558502 604894
rect 558586 604658 558822 604894
rect 558266 604338 558502 604574
rect 558586 604338 558822 604574
rect 558266 568658 558502 568894
rect 558586 568658 558822 568894
rect 558266 568338 558502 568574
rect 558586 568338 558822 568574
rect 558266 532658 558502 532894
rect 558586 532658 558822 532894
rect 558266 532338 558502 532574
rect 558586 532338 558822 532574
rect 558266 496658 558502 496894
rect 558586 496658 558822 496894
rect 558266 496338 558502 496574
rect 558586 496338 558822 496574
rect 558266 460658 558502 460894
rect 558586 460658 558822 460894
rect 558266 460338 558502 460574
rect 558586 460338 558822 460574
rect 558266 424658 558502 424894
rect 558586 424658 558822 424894
rect 558266 424338 558502 424574
rect 558586 424338 558822 424574
rect 558266 388658 558502 388894
rect 558586 388658 558822 388894
rect 558266 388338 558502 388574
rect 558586 388338 558822 388574
rect 558266 352658 558502 352894
rect 558586 352658 558822 352894
rect 558266 352338 558502 352574
rect 558586 352338 558822 352574
rect 558266 316658 558502 316894
rect 558586 316658 558822 316894
rect 558266 316338 558502 316574
rect 558586 316338 558822 316574
rect 558266 280658 558502 280894
rect 558586 280658 558822 280894
rect 558266 280338 558502 280574
rect 558586 280338 558822 280574
rect 558266 244658 558502 244894
rect 558586 244658 558822 244894
rect 558266 244338 558502 244574
rect 558586 244338 558822 244574
rect 558266 208658 558502 208894
rect 558586 208658 558822 208894
rect 558266 208338 558502 208574
rect 558586 208338 558822 208574
rect 558266 172658 558502 172894
rect 558586 172658 558822 172894
rect 558266 172338 558502 172574
rect 558586 172338 558822 172574
rect 558266 136658 558502 136894
rect 558586 136658 558822 136894
rect 558266 136338 558502 136574
rect 558586 136338 558822 136574
rect 558266 100658 558502 100894
rect 558586 100658 558822 100894
rect 558266 100338 558502 100574
rect 558586 100338 558822 100574
rect 558266 64658 558502 64894
rect 558586 64658 558822 64894
rect 558266 64338 558502 64574
rect 558586 64338 558822 64574
rect 558266 28658 558502 28894
rect 558586 28658 558822 28894
rect 558266 28338 558502 28574
rect 558586 28338 558822 28574
rect 560826 704602 561062 704838
rect 561146 704602 561382 704838
rect 560826 704282 561062 704518
rect 561146 704282 561382 704518
rect 560826 687218 561062 687454
rect 561146 687218 561382 687454
rect 560826 686898 561062 687134
rect 561146 686898 561382 687134
rect 560826 651218 561062 651454
rect 561146 651218 561382 651454
rect 560826 650898 561062 651134
rect 561146 650898 561382 651134
rect 560826 615218 561062 615454
rect 561146 615218 561382 615454
rect 560826 614898 561062 615134
rect 561146 614898 561382 615134
rect 560826 579218 561062 579454
rect 561146 579218 561382 579454
rect 560826 578898 561062 579134
rect 561146 578898 561382 579134
rect 560826 543218 561062 543454
rect 561146 543218 561382 543454
rect 560826 542898 561062 543134
rect 561146 542898 561382 543134
rect 560826 507218 561062 507454
rect 561146 507218 561382 507454
rect 560826 506898 561062 507134
rect 561146 506898 561382 507134
rect 560826 471218 561062 471454
rect 561146 471218 561382 471454
rect 560826 470898 561062 471134
rect 561146 470898 561382 471134
rect 560826 435218 561062 435454
rect 561146 435218 561382 435454
rect 560826 434898 561062 435134
rect 561146 434898 561382 435134
rect 560826 399218 561062 399454
rect 561146 399218 561382 399454
rect 560826 398898 561062 399134
rect 561146 398898 561382 399134
rect 560826 363218 561062 363454
rect 561146 363218 561382 363454
rect 560826 362898 561062 363134
rect 561146 362898 561382 363134
rect 560826 327218 561062 327454
rect 561146 327218 561382 327454
rect 560826 326898 561062 327134
rect 561146 326898 561382 327134
rect 560826 291218 561062 291454
rect 561146 291218 561382 291454
rect 560826 290898 561062 291134
rect 561146 290898 561382 291134
rect 560826 255218 561062 255454
rect 561146 255218 561382 255454
rect 560826 254898 561062 255134
rect 561146 254898 561382 255134
rect 560826 219218 561062 219454
rect 561146 219218 561382 219454
rect 560826 218898 561062 219134
rect 561146 218898 561382 219134
rect 560826 183218 561062 183454
rect 561146 183218 561382 183454
rect 560826 182898 561062 183134
rect 561146 182898 561382 183134
rect 560826 147218 561062 147454
rect 561146 147218 561382 147454
rect 560826 146898 561062 147134
rect 561146 146898 561382 147134
rect 560826 111218 561062 111454
rect 561146 111218 561382 111454
rect 560826 110898 561062 111134
rect 561146 110898 561382 111134
rect 560826 75218 561062 75454
rect 561146 75218 561382 75454
rect 560826 74898 561062 75134
rect 561146 74898 561382 75134
rect 560826 39218 561062 39454
rect 561146 39218 561382 39454
rect 560826 38898 561062 39134
rect 561146 38898 561382 39134
rect 560826 3218 561062 3454
rect 561146 3218 561382 3454
rect 560826 2898 561062 3134
rect 561146 2898 561382 3134
rect 560826 -582 561062 -346
rect 561146 -582 561382 -346
rect 560826 -902 561062 -666
rect 561146 -902 561382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 571986 710362 572222 710598
rect 572306 710362 572542 710598
rect 571986 710042 572222 710278
rect 572306 710042 572542 710278
rect 568266 708442 568502 708678
rect 568586 708442 568822 708678
rect 568266 708122 568502 708358
rect 568586 708122 568822 708358
rect 561986 680378 562222 680614
rect 562306 680378 562542 680614
rect 561986 680058 562222 680294
rect 562306 680058 562542 680294
rect 561986 644378 562222 644614
rect 562306 644378 562542 644614
rect 561986 644058 562222 644294
rect 562306 644058 562542 644294
rect 561986 608378 562222 608614
rect 562306 608378 562542 608614
rect 561986 608058 562222 608294
rect 562306 608058 562542 608294
rect 561986 572378 562222 572614
rect 562306 572378 562542 572614
rect 561986 572058 562222 572294
rect 562306 572058 562542 572294
rect 561986 536378 562222 536614
rect 562306 536378 562542 536614
rect 561986 536058 562222 536294
rect 562306 536058 562542 536294
rect 561986 500378 562222 500614
rect 562306 500378 562542 500614
rect 561986 500058 562222 500294
rect 562306 500058 562542 500294
rect 561986 464378 562222 464614
rect 562306 464378 562542 464614
rect 561986 464058 562222 464294
rect 562306 464058 562542 464294
rect 561986 428378 562222 428614
rect 562306 428378 562542 428614
rect 561986 428058 562222 428294
rect 562306 428058 562542 428294
rect 561986 392378 562222 392614
rect 562306 392378 562542 392614
rect 561986 392058 562222 392294
rect 562306 392058 562542 392294
rect 561986 356378 562222 356614
rect 562306 356378 562542 356614
rect 561986 356058 562222 356294
rect 562306 356058 562542 356294
rect 561986 320378 562222 320614
rect 562306 320378 562542 320614
rect 561986 320058 562222 320294
rect 562306 320058 562542 320294
rect 561986 284378 562222 284614
rect 562306 284378 562542 284614
rect 561986 284058 562222 284294
rect 562306 284058 562542 284294
rect 561986 248378 562222 248614
rect 562306 248378 562542 248614
rect 561986 248058 562222 248294
rect 562306 248058 562542 248294
rect 561986 212378 562222 212614
rect 562306 212378 562542 212614
rect 561986 212058 562222 212294
rect 562306 212058 562542 212294
rect 561986 176378 562222 176614
rect 562306 176378 562542 176614
rect 561986 176058 562222 176294
rect 562306 176058 562542 176294
rect 561986 140378 562222 140614
rect 562306 140378 562542 140614
rect 561986 140058 562222 140294
rect 562306 140058 562542 140294
rect 561986 104378 562222 104614
rect 562306 104378 562542 104614
rect 561986 104058 562222 104294
rect 562306 104058 562542 104294
rect 561986 68378 562222 68614
rect 562306 68378 562542 68614
rect 561986 68058 562222 68294
rect 562306 68058 562542 68294
rect 561986 32378 562222 32614
rect 562306 32378 562542 32614
rect 561986 32058 562222 32294
rect 562306 32058 562542 32294
rect 558266 -5382 558502 -5146
rect 558586 -5382 558822 -5146
rect 558266 -5702 558502 -5466
rect 558586 -5702 558822 -5466
rect 551986 -6342 552222 -6106
rect 552306 -6342 552542 -6106
rect 551986 -6662 552222 -6426
rect 552306 -6662 552542 -6426
rect 564546 706522 564782 706758
rect 564866 706522 565102 706758
rect 564546 706202 564782 706438
rect 564866 706202 565102 706438
rect 564546 690938 564782 691174
rect 564866 690938 565102 691174
rect 564546 690618 564782 690854
rect 564866 690618 565102 690854
rect 564546 654938 564782 655174
rect 564866 654938 565102 655174
rect 564546 654618 564782 654854
rect 564866 654618 565102 654854
rect 564546 618938 564782 619174
rect 564866 618938 565102 619174
rect 564546 618618 564782 618854
rect 564866 618618 565102 618854
rect 564546 582938 564782 583174
rect 564866 582938 565102 583174
rect 564546 582618 564782 582854
rect 564866 582618 565102 582854
rect 564546 546938 564782 547174
rect 564866 546938 565102 547174
rect 564546 546618 564782 546854
rect 564866 546618 565102 546854
rect 564546 510938 564782 511174
rect 564866 510938 565102 511174
rect 564546 510618 564782 510854
rect 564866 510618 565102 510854
rect 564546 474938 564782 475174
rect 564866 474938 565102 475174
rect 564546 474618 564782 474854
rect 564866 474618 565102 474854
rect 564546 438938 564782 439174
rect 564866 438938 565102 439174
rect 564546 438618 564782 438854
rect 564866 438618 565102 438854
rect 564546 402938 564782 403174
rect 564866 402938 565102 403174
rect 564546 402618 564782 402854
rect 564866 402618 565102 402854
rect 564546 366938 564782 367174
rect 564866 366938 565102 367174
rect 564546 366618 564782 366854
rect 564866 366618 565102 366854
rect 564546 330938 564782 331174
rect 564866 330938 565102 331174
rect 564546 330618 564782 330854
rect 564866 330618 565102 330854
rect 564546 294938 564782 295174
rect 564866 294938 565102 295174
rect 564546 294618 564782 294854
rect 564866 294618 565102 294854
rect 564546 258938 564782 259174
rect 564866 258938 565102 259174
rect 564546 258618 564782 258854
rect 564866 258618 565102 258854
rect 564546 222938 564782 223174
rect 564866 222938 565102 223174
rect 564546 222618 564782 222854
rect 564866 222618 565102 222854
rect 564546 186938 564782 187174
rect 564866 186938 565102 187174
rect 564546 186618 564782 186854
rect 564866 186618 565102 186854
rect 564546 150938 564782 151174
rect 564866 150938 565102 151174
rect 564546 150618 564782 150854
rect 564866 150618 565102 150854
rect 564546 114938 564782 115174
rect 564866 114938 565102 115174
rect 564546 114618 564782 114854
rect 564866 114618 565102 114854
rect 564546 78938 564782 79174
rect 564866 78938 565102 79174
rect 564546 78618 564782 78854
rect 564866 78618 565102 78854
rect 564546 42938 564782 43174
rect 564866 42938 565102 43174
rect 564546 42618 564782 42854
rect 564866 42618 565102 42854
rect 564546 6938 564782 7174
rect 564866 6938 565102 7174
rect 564546 6618 564782 6854
rect 564866 6618 565102 6854
rect 564546 -2502 564782 -2266
rect 564866 -2502 565102 -2266
rect 564546 -2822 564782 -2586
rect 564866 -2822 565102 -2586
rect 568266 694658 568502 694894
rect 568586 694658 568822 694894
rect 568266 694338 568502 694574
rect 568586 694338 568822 694574
rect 568266 658658 568502 658894
rect 568586 658658 568822 658894
rect 568266 658338 568502 658574
rect 568586 658338 568822 658574
rect 568266 622658 568502 622894
rect 568586 622658 568822 622894
rect 568266 622338 568502 622574
rect 568586 622338 568822 622574
rect 568266 586658 568502 586894
rect 568586 586658 568822 586894
rect 568266 586338 568502 586574
rect 568586 586338 568822 586574
rect 568266 550658 568502 550894
rect 568586 550658 568822 550894
rect 568266 550338 568502 550574
rect 568586 550338 568822 550574
rect 568266 514658 568502 514894
rect 568586 514658 568822 514894
rect 568266 514338 568502 514574
rect 568586 514338 568822 514574
rect 568266 478658 568502 478894
rect 568586 478658 568822 478894
rect 568266 478338 568502 478574
rect 568586 478338 568822 478574
rect 568266 442658 568502 442894
rect 568586 442658 568822 442894
rect 568266 442338 568502 442574
rect 568586 442338 568822 442574
rect 568266 406658 568502 406894
rect 568586 406658 568822 406894
rect 568266 406338 568502 406574
rect 568586 406338 568822 406574
rect 568266 370658 568502 370894
rect 568586 370658 568822 370894
rect 568266 370338 568502 370574
rect 568586 370338 568822 370574
rect 568266 334658 568502 334894
rect 568586 334658 568822 334894
rect 568266 334338 568502 334574
rect 568586 334338 568822 334574
rect 568266 298658 568502 298894
rect 568586 298658 568822 298894
rect 568266 298338 568502 298574
rect 568586 298338 568822 298574
rect 568266 262658 568502 262894
rect 568586 262658 568822 262894
rect 568266 262338 568502 262574
rect 568586 262338 568822 262574
rect 568266 226658 568502 226894
rect 568586 226658 568822 226894
rect 568266 226338 568502 226574
rect 568586 226338 568822 226574
rect 568266 190658 568502 190894
rect 568586 190658 568822 190894
rect 568266 190338 568502 190574
rect 568586 190338 568822 190574
rect 568266 154658 568502 154894
rect 568586 154658 568822 154894
rect 568266 154338 568502 154574
rect 568586 154338 568822 154574
rect 568266 118658 568502 118894
rect 568586 118658 568822 118894
rect 568266 118338 568502 118574
rect 568586 118338 568822 118574
rect 568266 82658 568502 82894
rect 568586 82658 568822 82894
rect 568266 82338 568502 82574
rect 568586 82338 568822 82574
rect 568266 46658 568502 46894
rect 568586 46658 568822 46894
rect 568266 46338 568502 46574
rect 568586 46338 568822 46574
rect 568266 10658 568502 10894
rect 568586 10658 568822 10894
rect 568266 10338 568502 10574
rect 568586 10338 568822 10574
rect 570826 705562 571062 705798
rect 571146 705562 571382 705798
rect 570826 705242 571062 705478
rect 571146 705242 571382 705478
rect 570826 669218 571062 669454
rect 571146 669218 571382 669454
rect 570826 668898 571062 669134
rect 571146 668898 571382 669134
rect 570826 633218 571062 633454
rect 571146 633218 571382 633454
rect 570826 632898 571062 633134
rect 571146 632898 571382 633134
rect 570826 597218 571062 597454
rect 571146 597218 571382 597454
rect 570826 596898 571062 597134
rect 571146 596898 571382 597134
rect 570826 561218 571062 561454
rect 571146 561218 571382 561454
rect 570826 560898 571062 561134
rect 571146 560898 571382 561134
rect 570826 525218 571062 525454
rect 571146 525218 571382 525454
rect 570826 524898 571062 525134
rect 571146 524898 571382 525134
rect 570826 489218 571062 489454
rect 571146 489218 571382 489454
rect 570826 488898 571062 489134
rect 571146 488898 571382 489134
rect 570826 453218 571062 453454
rect 571146 453218 571382 453454
rect 570826 452898 571062 453134
rect 571146 452898 571382 453134
rect 570826 417218 571062 417454
rect 571146 417218 571382 417454
rect 570826 416898 571062 417134
rect 571146 416898 571382 417134
rect 570826 381218 571062 381454
rect 571146 381218 571382 381454
rect 570826 380898 571062 381134
rect 571146 380898 571382 381134
rect 570826 345218 571062 345454
rect 571146 345218 571382 345454
rect 570826 344898 571062 345134
rect 571146 344898 571382 345134
rect 570826 309218 571062 309454
rect 571146 309218 571382 309454
rect 570826 308898 571062 309134
rect 571146 308898 571382 309134
rect 570826 273218 571062 273454
rect 571146 273218 571382 273454
rect 570826 272898 571062 273134
rect 571146 272898 571382 273134
rect 570826 237218 571062 237454
rect 571146 237218 571382 237454
rect 570826 236898 571062 237134
rect 571146 236898 571382 237134
rect 570826 201218 571062 201454
rect 571146 201218 571382 201454
rect 570826 200898 571062 201134
rect 571146 200898 571382 201134
rect 570826 165218 571062 165454
rect 571146 165218 571382 165454
rect 570826 164898 571062 165134
rect 571146 164898 571382 165134
rect 570826 129218 571062 129454
rect 571146 129218 571382 129454
rect 570826 128898 571062 129134
rect 571146 128898 571382 129134
rect 570826 93218 571062 93454
rect 571146 93218 571382 93454
rect 570826 92898 571062 93134
rect 571146 92898 571382 93134
rect 570826 57218 571062 57454
rect 571146 57218 571382 57454
rect 570826 56898 571062 57134
rect 571146 56898 571382 57134
rect 570826 21218 571062 21454
rect 571146 21218 571382 21454
rect 570826 20898 571062 21134
rect 571146 20898 571382 21134
rect 570826 -1542 571062 -1306
rect 571146 -1542 571382 -1306
rect 570826 -1862 571062 -1626
rect 571146 -1862 571382 -1626
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 578266 709402 578502 709638
rect 578586 709402 578822 709638
rect 578266 709082 578502 709318
rect 578586 709082 578822 709318
rect 571986 698378 572222 698614
rect 572306 698378 572542 698614
rect 571986 698058 572222 698294
rect 572306 698058 572542 698294
rect 571986 662378 572222 662614
rect 572306 662378 572542 662614
rect 571986 662058 572222 662294
rect 572306 662058 572542 662294
rect 571986 626378 572222 626614
rect 572306 626378 572542 626614
rect 571986 626058 572222 626294
rect 572306 626058 572542 626294
rect 571986 590378 572222 590614
rect 572306 590378 572542 590614
rect 571986 590058 572222 590294
rect 572306 590058 572542 590294
rect 571986 554378 572222 554614
rect 572306 554378 572542 554614
rect 571986 554058 572222 554294
rect 572306 554058 572542 554294
rect 571986 518378 572222 518614
rect 572306 518378 572542 518614
rect 571986 518058 572222 518294
rect 572306 518058 572542 518294
rect 571986 482378 572222 482614
rect 572306 482378 572542 482614
rect 571986 482058 572222 482294
rect 572306 482058 572542 482294
rect 571986 446378 572222 446614
rect 572306 446378 572542 446614
rect 571986 446058 572222 446294
rect 572306 446058 572542 446294
rect 571986 410378 572222 410614
rect 572306 410378 572542 410614
rect 571986 410058 572222 410294
rect 572306 410058 572542 410294
rect 571986 374378 572222 374614
rect 572306 374378 572542 374614
rect 571986 374058 572222 374294
rect 572306 374058 572542 374294
rect 571986 338378 572222 338614
rect 572306 338378 572542 338614
rect 571986 338058 572222 338294
rect 572306 338058 572542 338294
rect 571986 302378 572222 302614
rect 572306 302378 572542 302614
rect 571986 302058 572222 302294
rect 572306 302058 572542 302294
rect 571986 266378 572222 266614
rect 572306 266378 572542 266614
rect 571986 266058 572222 266294
rect 572306 266058 572542 266294
rect 571986 230378 572222 230614
rect 572306 230378 572542 230614
rect 571986 230058 572222 230294
rect 572306 230058 572542 230294
rect 571986 194378 572222 194614
rect 572306 194378 572542 194614
rect 571986 194058 572222 194294
rect 572306 194058 572542 194294
rect 571986 158378 572222 158614
rect 572306 158378 572542 158614
rect 571986 158058 572222 158294
rect 572306 158058 572542 158294
rect 571986 122378 572222 122614
rect 572306 122378 572542 122614
rect 571986 122058 572222 122294
rect 572306 122058 572542 122294
rect 571986 86378 572222 86614
rect 572306 86378 572542 86614
rect 571986 86058 572222 86294
rect 572306 86058 572542 86294
rect 571986 50378 572222 50614
rect 572306 50378 572542 50614
rect 571986 50058 572222 50294
rect 572306 50058 572542 50294
rect 571986 14378 572222 14614
rect 572306 14378 572542 14614
rect 571986 14058 572222 14294
rect 572306 14058 572542 14294
rect 568266 -4422 568502 -4186
rect 568586 -4422 568822 -4186
rect 568266 -4742 568502 -4506
rect 568586 -4742 568822 -4506
rect 561986 -7302 562222 -7066
rect 562306 -7302 562542 -7066
rect 561986 -7622 562222 -7386
rect 562306 -7622 562542 -7386
rect 574546 707482 574782 707718
rect 574866 707482 575102 707718
rect 574546 707162 574782 707398
rect 574866 707162 575102 707398
rect 574546 672938 574782 673174
rect 574866 672938 575102 673174
rect 574546 672618 574782 672854
rect 574866 672618 575102 672854
rect 574546 636938 574782 637174
rect 574866 636938 575102 637174
rect 574546 636618 574782 636854
rect 574866 636618 575102 636854
rect 574546 600938 574782 601174
rect 574866 600938 575102 601174
rect 574546 600618 574782 600854
rect 574866 600618 575102 600854
rect 574546 564938 574782 565174
rect 574866 564938 575102 565174
rect 574546 564618 574782 564854
rect 574866 564618 575102 564854
rect 574546 528938 574782 529174
rect 574866 528938 575102 529174
rect 574546 528618 574782 528854
rect 574866 528618 575102 528854
rect 574546 492938 574782 493174
rect 574866 492938 575102 493174
rect 574546 492618 574782 492854
rect 574866 492618 575102 492854
rect 574546 456938 574782 457174
rect 574866 456938 575102 457174
rect 574546 456618 574782 456854
rect 574866 456618 575102 456854
rect 574546 420938 574782 421174
rect 574866 420938 575102 421174
rect 574546 420618 574782 420854
rect 574866 420618 575102 420854
rect 574546 384938 574782 385174
rect 574866 384938 575102 385174
rect 574546 384618 574782 384854
rect 574866 384618 575102 384854
rect 574546 348938 574782 349174
rect 574866 348938 575102 349174
rect 574546 348618 574782 348854
rect 574866 348618 575102 348854
rect 574546 312938 574782 313174
rect 574866 312938 575102 313174
rect 574546 312618 574782 312854
rect 574866 312618 575102 312854
rect 574546 276938 574782 277174
rect 574866 276938 575102 277174
rect 574546 276618 574782 276854
rect 574866 276618 575102 276854
rect 574546 240938 574782 241174
rect 574866 240938 575102 241174
rect 574546 240618 574782 240854
rect 574866 240618 575102 240854
rect 574546 204938 574782 205174
rect 574866 204938 575102 205174
rect 574546 204618 574782 204854
rect 574866 204618 575102 204854
rect 574546 168938 574782 169174
rect 574866 168938 575102 169174
rect 574546 168618 574782 168854
rect 574866 168618 575102 168854
rect 574546 132938 574782 133174
rect 574866 132938 575102 133174
rect 574546 132618 574782 132854
rect 574866 132618 575102 132854
rect 574546 96938 574782 97174
rect 574866 96938 575102 97174
rect 574546 96618 574782 96854
rect 574866 96618 575102 96854
rect 574546 60938 574782 61174
rect 574866 60938 575102 61174
rect 574546 60618 574782 60854
rect 574866 60618 575102 60854
rect 574546 24938 574782 25174
rect 574866 24938 575102 25174
rect 574546 24618 574782 24854
rect 574866 24618 575102 24854
rect 574546 -3462 574782 -3226
rect 574866 -3462 575102 -3226
rect 574546 -3782 574782 -3546
rect 574866 -3782 575102 -3546
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 578266 676658 578502 676894
rect 578586 676658 578822 676894
rect 578266 676338 578502 676574
rect 578586 676338 578822 676574
rect 578266 640658 578502 640894
rect 578586 640658 578822 640894
rect 578266 640338 578502 640574
rect 578586 640338 578822 640574
rect 578266 604658 578502 604894
rect 578586 604658 578822 604894
rect 578266 604338 578502 604574
rect 578586 604338 578822 604574
rect 578266 568658 578502 568894
rect 578586 568658 578822 568894
rect 578266 568338 578502 568574
rect 578586 568338 578822 568574
rect 578266 532658 578502 532894
rect 578586 532658 578822 532894
rect 578266 532338 578502 532574
rect 578586 532338 578822 532574
rect 578266 496658 578502 496894
rect 578586 496658 578822 496894
rect 578266 496338 578502 496574
rect 578586 496338 578822 496574
rect 578266 460658 578502 460894
rect 578586 460658 578822 460894
rect 578266 460338 578502 460574
rect 578586 460338 578822 460574
rect 578266 424658 578502 424894
rect 578586 424658 578822 424894
rect 578266 424338 578502 424574
rect 578586 424338 578822 424574
rect 578266 388658 578502 388894
rect 578586 388658 578822 388894
rect 578266 388338 578502 388574
rect 578586 388338 578822 388574
rect 578266 352658 578502 352894
rect 578586 352658 578822 352894
rect 578266 352338 578502 352574
rect 578586 352338 578822 352574
rect 578266 316658 578502 316894
rect 578586 316658 578822 316894
rect 578266 316338 578502 316574
rect 578586 316338 578822 316574
rect 578266 280658 578502 280894
rect 578586 280658 578822 280894
rect 578266 280338 578502 280574
rect 578586 280338 578822 280574
rect 578266 244658 578502 244894
rect 578586 244658 578822 244894
rect 578266 244338 578502 244574
rect 578586 244338 578822 244574
rect 578266 208658 578502 208894
rect 578586 208658 578822 208894
rect 578266 208338 578502 208574
rect 578586 208338 578822 208574
rect 578266 172658 578502 172894
rect 578586 172658 578822 172894
rect 578266 172338 578502 172574
rect 578586 172338 578822 172574
rect 578266 136658 578502 136894
rect 578586 136658 578822 136894
rect 578266 136338 578502 136574
rect 578586 136338 578822 136574
rect 578266 100658 578502 100894
rect 578586 100658 578822 100894
rect 578266 100338 578502 100574
rect 578586 100338 578822 100574
rect 578266 64658 578502 64894
rect 578586 64658 578822 64894
rect 578266 64338 578502 64574
rect 578586 64338 578822 64574
rect 578266 28658 578502 28894
rect 578586 28658 578822 28894
rect 578266 28338 578502 28574
rect 578586 28338 578822 28574
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 580826 704602 581062 704838
rect 581146 704602 581382 704838
rect 580826 704282 581062 704518
rect 581146 704282 581382 704518
rect 580826 687218 581062 687454
rect 581146 687218 581382 687454
rect 580826 686898 581062 687134
rect 581146 686898 581382 687134
rect 580826 651218 581062 651454
rect 581146 651218 581382 651454
rect 580826 650898 581062 651134
rect 581146 650898 581382 651134
rect 580826 615218 581062 615454
rect 581146 615218 581382 615454
rect 580826 614898 581062 615134
rect 581146 614898 581382 615134
rect 580826 579218 581062 579454
rect 581146 579218 581382 579454
rect 580826 578898 581062 579134
rect 581146 578898 581382 579134
rect 580826 543218 581062 543454
rect 581146 543218 581382 543454
rect 580826 542898 581062 543134
rect 581146 542898 581382 543134
rect 580826 507218 581062 507454
rect 581146 507218 581382 507454
rect 580826 506898 581062 507134
rect 581146 506898 581382 507134
rect 580826 471218 581062 471454
rect 581146 471218 581382 471454
rect 580826 470898 581062 471134
rect 581146 470898 581382 471134
rect 580826 435218 581062 435454
rect 581146 435218 581382 435454
rect 580826 434898 581062 435134
rect 581146 434898 581382 435134
rect 580826 399218 581062 399454
rect 581146 399218 581382 399454
rect 580826 398898 581062 399134
rect 581146 398898 581382 399134
rect 580826 363218 581062 363454
rect 581146 363218 581382 363454
rect 580826 362898 581062 363134
rect 581146 362898 581382 363134
rect 580826 327218 581062 327454
rect 581146 327218 581382 327454
rect 580826 326898 581062 327134
rect 581146 326898 581382 327134
rect 580826 291218 581062 291454
rect 581146 291218 581382 291454
rect 580826 290898 581062 291134
rect 581146 290898 581382 291134
rect 580826 255218 581062 255454
rect 581146 255218 581382 255454
rect 580826 254898 581062 255134
rect 581146 254898 581382 255134
rect 580826 219218 581062 219454
rect 581146 219218 581382 219454
rect 580826 218898 581062 219134
rect 581146 218898 581382 219134
rect 580826 183218 581062 183454
rect 581146 183218 581382 183454
rect 580826 182898 581062 183134
rect 581146 182898 581382 183134
rect 580826 147218 581062 147454
rect 581146 147218 581382 147454
rect 580826 146898 581062 147134
rect 581146 146898 581382 147134
rect 580826 111218 581062 111454
rect 581146 111218 581382 111454
rect 580826 110898 581062 111134
rect 581146 110898 581382 111134
rect 580826 75218 581062 75454
rect 581146 75218 581382 75454
rect 580826 74898 581062 75134
rect 581146 74898 581382 75134
rect 580826 39218 581062 39454
rect 581146 39218 581382 39454
rect 580826 38898 581062 39134
rect 581146 38898 581382 39134
rect 580826 3218 581062 3454
rect 581146 3218 581382 3454
rect 580826 2898 581062 3134
rect 581146 2898 581382 3134
rect 580826 -582 581062 -346
rect 581146 -582 581382 -346
rect 580826 -902 581062 -666
rect 581146 -902 581382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 578266 -5382 578502 -5146
rect 578586 -5382 578822 -5146
rect 578266 -5702 578502 -5466
rect 578586 -5702 578822 -5466
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 571986 -6342 572222 -6106
rect 572306 -6342 572542 -6106
rect 571986 -6662 572222 -6426
rect 572306 -6662 572542 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 21986 711558
rect 22222 711322 22306 711558
rect 22542 711322 41986 711558
rect 42222 711322 42306 711558
rect 42542 711322 61986 711558
rect 62222 711322 62306 711558
rect 62542 711322 81986 711558
rect 82222 711322 82306 711558
rect 82542 711322 101986 711558
rect 102222 711322 102306 711558
rect 102542 711322 121986 711558
rect 122222 711322 122306 711558
rect 122542 711322 141986 711558
rect 142222 711322 142306 711558
rect 142542 711322 161986 711558
rect 162222 711322 162306 711558
rect 162542 711322 181986 711558
rect 182222 711322 182306 711558
rect 182542 711322 201986 711558
rect 202222 711322 202306 711558
rect 202542 711322 221986 711558
rect 222222 711322 222306 711558
rect 222542 711322 241986 711558
rect 242222 711322 242306 711558
rect 242542 711322 261986 711558
rect 262222 711322 262306 711558
rect 262542 711322 281986 711558
rect 282222 711322 282306 711558
rect 282542 711322 301986 711558
rect 302222 711322 302306 711558
rect 302542 711322 321986 711558
rect 322222 711322 322306 711558
rect 322542 711322 341986 711558
rect 342222 711322 342306 711558
rect 342542 711322 361986 711558
rect 362222 711322 362306 711558
rect 362542 711322 381986 711558
rect 382222 711322 382306 711558
rect 382542 711322 401986 711558
rect 402222 711322 402306 711558
rect 402542 711322 421986 711558
rect 422222 711322 422306 711558
rect 422542 711322 441986 711558
rect 442222 711322 442306 711558
rect 442542 711322 461986 711558
rect 462222 711322 462306 711558
rect 462542 711322 481986 711558
rect 482222 711322 482306 711558
rect 482542 711322 501986 711558
rect 502222 711322 502306 711558
rect 502542 711322 521986 711558
rect 522222 711322 522306 711558
rect 522542 711322 541986 711558
rect 542222 711322 542306 711558
rect 542542 711322 561986 711558
rect 562222 711322 562306 711558
rect 562542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 21986 711238
rect 22222 711002 22306 711238
rect 22542 711002 41986 711238
rect 42222 711002 42306 711238
rect 42542 711002 61986 711238
rect 62222 711002 62306 711238
rect 62542 711002 81986 711238
rect 82222 711002 82306 711238
rect 82542 711002 101986 711238
rect 102222 711002 102306 711238
rect 102542 711002 121986 711238
rect 122222 711002 122306 711238
rect 122542 711002 141986 711238
rect 142222 711002 142306 711238
rect 142542 711002 161986 711238
rect 162222 711002 162306 711238
rect 162542 711002 181986 711238
rect 182222 711002 182306 711238
rect 182542 711002 201986 711238
rect 202222 711002 202306 711238
rect 202542 711002 221986 711238
rect 222222 711002 222306 711238
rect 222542 711002 241986 711238
rect 242222 711002 242306 711238
rect 242542 711002 261986 711238
rect 262222 711002 262306 711238
rect 262542 711002 281986 711238
rect 282222 711002 282306 711238
rect 282542 711002 301986 711238
rect 302222 711002 302306 711238
rect 302542 711002 321986 711238
rect 322222 711002 322306 711238
rect 322542 711002 341986 711238
rect 342222 711002 342306 711238
rect 342542 711002 361986 711238
rect 362222 711002 362306 711238
rect 362542 711002 381986 711238
rect 382222 711002 382306 711238
rect 382542 711002 401986 711238
rect 402222 711002 402306 711238
rect 402542 711002 421986 711238
rect 422222 711002 422306 711238
rect 422542 711002 441986 711238
rect 442222 711002 442306 711238
rect 442542 711002 461986 711238
rect 462222 711002 462306 711238
rect 462542 711002 481986 711238
rect 482222 711002 482306 711238
rect 482542 711002 501986 711238
rect 502222 711002 502306 711238
rect 502542 711002 521986 711238
rect 522222 711002 522306 711238
rect 522542 711002 541986 711238
rect 542222 711002 542306 711238
rect 542542 711002 561986 711238
rect 562222 711002 562306 711238
rect 562542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 11986 710598
rect 12222 710362 12306 710598
rect 12542 710362 31986 710598
rect 32222 710362 32306 710598
rect 32542 710362 51986 710598
rect 52222 710362 52306 710598
rect 52542 710362 71986 710598
rect 72222 710362 72306 710598
rect 72542 710362 91986 710598
rect 92222 710362 92306 710598
rect 92542 710362 111986 710598
rect 112222 710362 112306 710598
rect 112542 710362 131986 710598
rect 132222 710362 132306 710598
rect 132542 710362 151986 710598
rect 152222 710362 152306 710598
rect 152542 710362 171986 710598
rect 172222 710362 172306 710598
rect 172542 710362 191986 710598
rect 192222 710362 192306 710598
rect 192542 710362 211986 710598
rect 212222 710362 212306 710598
rect 212542 710362 231986 710598
rect 232222 710362 232306 710598
rect 232542 710362 251986 710598
rect 252222 710362 252306 710598
rect 252542 710362 271986 710598
rect 272222 710362 272306 710598
rect 272542 710362 291986 710598
rect 292222 710362 292306 710598
rect 292542 710362 311986 710598
rect 312222 710362 312306 710598
rect 312542 710362 331986 710598
rect 332222 710362 332306 710598
rect 332542 710362 351986 710598
rect 352222 710362 352306 710598
rect 352542 710362 371986 710598
rect 372222 710362 372306 710598
rect 372542 710362 391986 710598
rect 392222 710362 392306 710598
rect 392542 710362 411986 710598
rect 412222 710362 412306 710598
rect 412542 710362 431986 710598
rect 432222 710362 432306 710598
rect 432542 710362 451986 710598
rect 452222 710362 452306 710598
rect 452542 710362 471986 710598
rect 472222 710362 472306 710598
rect 472542 710362 491986 710598
rect 492222 710362 492306 710598
rect 492542 710362 511986 710598
rect 512222 710362 512306 710598
rect 512542 710362 531986 710598
rect 532222 710362 532306 710598
rect 532542 710362 551986 710598
rect 552222 710362 552306 710598
rect 552542 710362 571986 710598
rect 572222 710362 572306 710598
rect 572542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 11986 710278
rect 12222 710042 12306 710278
rect 12542 710042 31986 710278
rect 32222 710042 32306 710278
rect 32542 710042 51986 710278
rect 52222 710042 52306 710278
rect 52542 710042 71986 710278
rect 72222 710042 72306 710278
rect 72542 710042 91986 710278
rect 92222 710042 92306 710278
rect 92542 710042 111986 710278
rect 112222 710042 112306 710278
rect 112542 710042 131986 710278
rect 132222 710042 132306 710278
rect 132542 710042 151986 710278
rect 152222 710042 152306 710278
rect 152542 710042 171986 710278
rect 172222 710042 172306 710278
rect 172542 710042 191986 710278
rect 192222 710042 192306 710278
rect 192542 710042 211986 710278
rect 212222 710042 212306 710278
rect 212542 710042 231986 710278
rect 232222 710042 232306 710278
rect 232542 710042 251986 710278
rect 252222 710042 252306 710278
rect 252542 710042 271986 710278
rect 272222 710042 272306 710278
rect 272542 710042 291986 710278
rect 292222 710042 292306 710278
rect 292542 710042 311986 710278
rect 312222 710042 312306 710278
rect 312542 710042 331986 710278
rect 332222 710042 332306 710278
rect 332542 710042 351986 710278
rect 352222 710042 352306 710278
rect 352542 710042 371986 710278
rect 372222 710042 372306 710278
rect 372542 710042 391986 710278
rect 392222 710042 392306 710278
rect 392542 710042 411986 710278
rect 412222 710042 412306 710278
rect 412542 710042 431986 710278
rect 432222 710042 432306 710278
rect 432542 710042 451986 710278
rect 452222 710042 452306 710278
rect 452542 710042 471986 710278
rect 472222 710042 472306 710278
rect 472542 710042 491986 710278
rect 492222 710042 492306 710278
rect 492542 710042 511986 710278
rect 512222 710042 512306 710278
rect 512542 710042 531986 710278
rect 532222 710042 532306 710278
rect 532542 710042 551986 710278
rect 552222 710042 552306 710278
rect 552542 710042 571986 710278
rect 572222 710042 572306 710278
rect 572542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 18266 709638
rect 18502 709402 18586 709638
rect 18822 709402 38266 709638
rect 38502 709402 38586 709638
rect 38822 709402 58266 709638
rect 58502 709402 58586 709638
rect 58822 709402 78266 709638
rect 78502 709402 78586 709638
rect 78822 709402 98266 709638
rect 98502 709402 98586 709638
rect 98822 709402 118266 709638
rect 118502 709402 118586 709638
rect 118822 709402 138266 709638
rect 138502 709402 138586 709638
rect 138822 709402 158266 709638
rect 158502 709402 158586 709638
rect 158822 709402 178266 709638
rect 178502 709402 178586 709638
rect 178822 709402 198266 709638
rect 198502 709402 198586 709638
rect 198822 709402 218266 709638
rect 218502 709402 218586 709638
rect 218822 709402 238266 709638
rect 238502 709402 238586 709638
rect 238822 709402 258266 709638
rect 258502 709402 258586 709638
rect 258822 709402 278266 709638
rect 278502 709402 278586 709638
rect 278822 709402 298266 709638
rect 298502 709402 298586 709638
rect 298822 709402 318266 709638
rect 318502 709402 318586 709638
rect 318822 709402 338266 709638
rect 338502 709402 338586 709638
rect 338822 709402 358266 709638
rect 358502 709402 358586 709638
rect 358822 709402 378266 709638
rect 378502 709402 378586 709638
rect 378822 709402 398266 709638
rect 398502 709402 398586 709638
rect 398822 709402 418266 709638
rect 418502 709402 418586 709638
rect 418822 709402 438266 709638
rect 438502 709402 438586 709638
rect 438822 709402 458266 709638
rect 458502 709402 458586 709638
rect 458822 709402 478266 709638
rect 478502 709402 478586 709638
rect 478822 709402 498266 709638
rect 498502 709402 498586 709638
rect 498822 709402 518266 709638
rect 518502 709402 518586 709638
rect 518822 709402 538266 709638
rect 538502 709402 538586 709638
rect 538822 709402 558266 709638
rect 558502 709402 558586 709638
rect 558822 709402 578266 709638
rect 578502 709402 578586 709638
rect 578822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 18266 709318
rect 18502 709082 18586 709318
rect 18822 709082 38266 709318
rect 38502 709082 38586 709318
rect 38822 709082 58266 709318
rect 58502 709082 58586 709318
rect 58822 709082 78266 709318
rect 78502 709082 78586 709318
rect 78822 709082 98266 709318
rect 98502 709082 98586 709318
rect 98822 709082 118266 709318
rect 118502 709082 118586 709318
rect 118822 709082 138266 709318
rect 138502 709082 138586 709318
rect 138822 709082 158266 709318
rect 158502 709082 158586 709318
rect 158822 709082 178266 709318
rect 178502 709082 178586 709318
rect 178822 709082 198266 709318
rect 198502 709082 198586 709318
rect 198822 709082 218266 709318
rect 218502 709082 218586 709318
rect 218822 709082 238266 709318
rect 238502 709082 238586 709318
rect 238822 709082 258266 709318
rect 258502 709082 258586 709318
rect 258822 709082 278266 709318
rect 278502 709082 278586 709318
rect 278822 709082 298266 709318
rect 298502 709082 298586 709318
rect 298822 709082 318266 709318
rect 318502 709082 318586 709318
rect 318822 709082 338266 709318
rect 338502 709082 338586 709318
rect 338822 709082 358266 709318
rect 358502 709082 358586 709318
rect 358822 709082 378266 709318
rect 378502 709082 378586 709318
rect 378822 709082 398266 709318
rect 398502 709082 398586 709318
rect 398822 709082 418266 709318
rect 418502 709082 418586 709318
rect 418822 709082 438266 709318
rect 438502 709082 438586 709318
rect 438822 709082 458266 709318
rect 458502 709082 458586 709318
rect 458822 709082 478266 709318
rect 478502 709082 478586 709318
rect 478822 709082 498266 709318
rect 498502 709082 498586 709318
rect 498822 709082 518266 709318
rect 518502 709082 518586 709318
rect 518822 709082 538266 709318
rect 538502 709082 538586 709318
rect 538822 709082 558266 709318
rect 558502 709082 558586 709318
rect 558822 709082 578266 709318
rect 578502 709082 578586 709318
rect 578822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 8266 708678
rect 8502 708442 8586 708678
rect 8822 708442 28266 708678
rect 28502 708442 28586 708678
rect 28822 708442 48266 708678
rect 48502 708442 48586 708678
rect 48822 708442 68266 708678
rect 68502 708442 68586 708678
rect 68822 708442 88266 708678
rect 88502 708442 88586 708678
rect 88822 708442 108266 708678
rect 108502 708442 108586 708678
rect 108822 708442 128266 708678
rect 128502 708442 128586 708678
rect 128822 708442 148266 708678
rect 148502 708442 148586 708678
rect 148822 708442 168266 708678
rect 168502 708442 168586 708678
rect 168822 708442 188266 708678
rect 188502 708442 188586 708678
rect 188822 708442 208266 708678
rect 208502 708442 208586 708678
rect 208822 708442 228266 708678
rect 228502 708442 228586 708678
rect 228822 708442 248266 708678
rect 248502 708442 248586 708678
rect 248822 708442 268266 708678
rect 268502 708442 268586 708678
rect 268822 708442 288266 708678
rect 288502 708442 288586 708678
rect 288822 708442 308266 708678
rect 308502 708442 308586 708678
rect 308822 708442 328266 708678
rect 328502 708442 328586 708678
rect 328822 708442 348266 708678
rect 348502 708442 348586 708678
rect 348822 708442 368266 708678
rect 368502 708442 368586 708678
rect 368822 708442 388266 708678
rect 388502 708442 388586 708678
rect 388822 708442 408266 708678
rect 408502 708442 408586 708678
rect 408822 708442 428266 708678
rect 428502 708442 428586 708678
rect 428822 708442 448266 708678
rect 448502 708442 448586 708678
rect 448822 708442 468266 708678
rect 468502 708442 468586 708678
rect 468822 708442 488266 708678
rect 488502 708442 488586 708678
rect 488822 708442 508266 708678
rect 508502 708442 508586 708678
rect 508822 708442 528266 708678
rect 528502 708442 528586 708678
rect 528822 708442 548266 708678
rect 548502 708442 548586 708678
rect 548822 708442 568266 708678
rect 568502 708442 568586 708678
rect 568822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 8266 708358
rect 8502 708122 8586 708358
rect 8822 708122 28266 708358
rect 28502 708122 28586 708358
rect 28822 708122 48266 708358
rect 48502 708122 48586 708358
rect 48822 708122 68266 708358
rect 68502 708122 68586 708358
rect 68822 708122 88266 708358
rect 88502 708122 88586 708358
rect 88822 708122 108266 708358
rect 108502 708122 108586 708358
rect 108822 708122 128266 708358
rect 128502 708122 128586 708358
rect 128822 708122 148266 708358
rect 148502 708122 148586 708358
rect 148822 708122 168266 708358
rect 168502 708122 168586 708358
rect 168822 708122 188266 708358
rect 188502 708122 188586 708358
rect 188822 708122 208266 708358
rect 208502 708122 208586 708358
rect 208822 708122 228266 708358
rect 228502 708122 228586 708358
rect 228822 708122 248266 708358
rect 248502 708122 248586 708358
rect 248822 708122 268266 708358
rect 268502 708122 268586 708358
rect 268822 708122 288266 708358
rect 288502 708122 288586 708358
rect 288822 708122 308266 708358
rect 308502 708122 308586 708358
rect 308822 708122 328266 708358
rect 328502 708122 328586 708358
rect 328822 708122 348266 708358
rect 348502 708122 348586 708358
rect 348822 708122 368266 708358
rect 368502 708122 368586 708358
rect 368822 708122 388266 708358
rect 388502 708122 388586 708358
rect 388822 708122 408266 708358
rect 408502 708122 408586 708358
rect 408822 708122 428266 708358
rect 428502 708122 428586 708358
rect 428822 708122 448266 708358
rect 448502 708122 448586 708358
rect 448822 708122 468266 708358
rect 468502 708122 468586 708358
rect 468822 708122 488266 708358
rect 488502 708122 488586 708358
rect 488822 708122 508266 708358
rect 508502 708122 508586 708358
rect 508822 708122 528266 708358
rect 528502 708122 528586 708358
rect 528822 708122 548266 708358
rect 548502 708122 548586 708358
rect 548822 708122 568266 708358
rect 568502 708122 568586 708358
rect 568822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 14546 707718
rect 14782 707482 14866 707718
rect 15102 707482 34546 707718
rect 34782 707482 34866 707718
rect 35102 707482 54546 707718
rect 54782 707482 54866 707718
rect 55102 707482 74546 707718
rect 74782 707482 74866 707718
rect 75102 707482 94546 707718
rect 94782 707482 94866 707718
rect 95102 707482 114546 707718
rect 114782 707482 114866 707718
rect 115102 707482 134546 707718
rect 134782 707482 134866 707718
rect 135102 707482 154546 707718
rect 154782 707482 154866 707718
rect 155102 707482 174546 707718
rect 174782 707482 174866 707718
rect 175102 707482 194546 707718
rect 194782 707482 194866 707718
rect 195102 707482 214546 707718
rect 214782 707482 214866 707718
rect 215102 707482 234546 707718
rect 234782 707482 234866 707718
rect 235102 707482 254546 707718
rect 254782 707482 254866 707718
rect 255102 707482 274546 707718
rect 274782 707482 274866 707718
rect 275102 707482 294546 707718
rect 294782 707482 294866 707718
rect 295102 707482 314546 707718
rect 314782 707482 314866 707718
rect 315102 707482 334546 707718
rect 334782 707482 334866 707718
rect 335102 707482 354546 707718
rect 354782 707482 354866 707718
rect 355102 707482 374546 707718
rect 374782 707482 374866 707718
rect 375102 707482 394546 707718
rect 394782 707482 394866 707718
rect 395102 707482 414546 707718
rect 414782 707482 414866 707718
rect 415102 707482 434546 707718
rect 434782 707482 434866 707718
rect 435102 707482 454546 707718
rect 454782 707482 454866 707718
rect 455102 707482 474546 707718
rect 474782 707482 474866 707718
rect 475102 707482 494546 707718
rect 494782 707482 494866 707718
rect 495102 707482 514546 707718
rect 514782 707482 514866 707718
rect 515102 707482 534546 707718
rect 534782 707482 534866 707718
rect 535102 707482 554546 707718
rect 554782 707482 554866 707718
rect 555102 707482 574546 707718
rect 574782 707482 574866 707718
rect 575102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 14546 707398
rect 14782 707162 14866 707398
rect 15102 707162 34546 707398
rect 34782 707162 34866 707398
rect 35102 707162 54546 707398
rect 54782 707162 54866 707398
rect 55102 707162 74546 707398
rect 74782 707162 74866 707398
rect 75102 707162 94546 707398
rect 94782 707162 94866 707398
rect 95102 707162 114546 707398
rect 114782 707162 114866 707398
rect 115102 707162 134546 707398
rect 134782 707162 134866 707398
rect 135102 707162 154546 707398
rect 154782 707162 154866 707398
rect 155102 707162 174546 707398
rect 174782 707162 174866 707398
rect 175102 707162 194546 707398
rect 194782 707162 194866 707398
rect 195102 707162 214546 707398
rect 214782 707162 214866 707398
rect 215102 707162 234546 707398
rect 234782 707162 234866 707398
rect 235102 707162 254546 707398
rect 254782 707162 254866 707398
rect 255102 707162 274546 707398
rect 274782 707162 274866 707398
rect 275102 707162 294546 707398
rect 294782 707162 294866 707398
rect 295102 707162 314546 707398
rect 314782 707162 314866 707398
rect 315102 707162 334546 707398
rect 334782 707162 334866 707398
rect 335102 707162 354546 707398
rect 354782 707162 354866 707398
rect 355102 707162 374546 707398
rect 374782 707162 374866 707398
rect 375102 707162 394546 707398
rect 394782 707162 394866 707398
rect 395102 707162 414546 707398
rect 414782 707162 414866 707398
rect 415102 707162 434546 707398
rect 434782 707162 434866 707398
rect 435102 707162 454546 707398
rect 454782 707162 454866 707398
rect 455102 707162 474546 707398
rect 474782 707162 474866 707398
rect 475102 707162 494546 707398
rect 494782 707162 494866 707398
rect 495102 707162 514546 707398
rect 514782 707162 514866 707398
rect 515102 707162 534546 707398
rect 534782 707162 534866 707398
rect 535102 707162 554546 707398
rect 554782 707162 554866 707398
rect 555102 707162 574546 707398
rect 574782 707162 574866 707398
rect 575102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 4546 706758
rect 4782 706522 4866 706758
rect 5102 706522 24546 706758
rect 24782 706522 24866 706758
rect 25102 706522 44546 706758
rect 44782 706522 44866 706758
rect 45102 706522 64546 706758
rect 64782 706522 64866 706758
rect 65102 706522 84546 706758
rect 84782 706522 84866 706758
rect 85102 706522 104546 706758
rect 104782 706522 104866 706758
rect 105102 706522 124546 706758
rect 124782 706522 124866 706758
rect 125102 706522 144546 706758
rect 144782 706522 144866 706758
rect 145102 706522 164546 706758
rect 164782 706522 164866 706758
rect 165102 706522 184546 706758
rect 184782 706522 184866 706758
rect 185102 706522 204546 706758
rect 204782 706522 204866 706758
rect 205102 706522 224546 706758
rect 224782 706522 224866 706758
rect 225102 706522 244546 706758
rect 244782 706522 244866 706758
rect 245102 706522 264546 706758
rect 264782 706522 264866 706758
rect 265102 706522 284546 706758
rect 284782 706522 284866 706758
rect 285102 706522 304546 706758
rect 304782 706522 304866 706758
rect 305102 706522 324546 706758
rect 324782 706522 324866 706758
rect 325102 706522 344546 706758
rect 344782 706522 344866 706758
rect 345102 706522 364546 706758
rect 364782 706522 364866 706758
rect 365102 706522 384546 706758
rect 384782 706522 384866 706758
rect 385102 706522 404546 706758
rect 404782 706522 404866 706758
rect 405102 706522 424546 706758
rect 424782 706522 424866 706758
rect 425102 706522 444546 706758
rect 444782 706522 444866 706758
rect 445102 706522 464546 706758
rect 464782 706522 464866 706758
rect 465102 706522 484546 706758
rect 484782 706522 484866 706758
rect 485102 706522 504546 706758
rect 504782 706522 504866 706758
rect 505102 706522 524546 706758
rect 524782 706522 524866 706758
rect 525102 706522 544546 706758
rect 544782 706522 544866 706758
rect 545102 706522 564546 706758
rect 564782 706522 564866 706758
rect 565102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 4546 706438
rect 4782 706202 4866 706438
rect 5102 706202 24546 706438
rect 24782 706202 24866 706438
rect 25102 706202 44546 706438
rect 44782 706202 44866 706438
rect 45102 706202 64546 706438
rect 64782 706202 64866 706438
rect 65102 706202 84546 706438
rect 84782 706202 84866 706438
rect 85102 706202 104546 706438
rect 104782 706202 104866 706438
rect 105102 706202 124546 706438
rect 124782 706202 124866 706438
rect 125102 706202 144546 706438
rect 144782 706202 144866 706438
rect 145102 706202 164546 706438
rect 164782 706202 164866 706438
rect 165102 706202 184546 706438
rect 184782 706202 184866 706438
rect 185102 706202 204546 706438
rect 204782 706202 204866 706438
rect 205102 706202 224546 706438
rect 224782 706202 224866 706438
rect 225102 706202 244546 706438
rect 244782 706202 244866 706438
rect 245102 706202 264546 706438
rect 264782 706202 264866 706438
rect 265102 706202 284546 706438
rect 284782 706202 284866 706438
rect 285102 706202 304546 706438
rect 304782 706202 304866 706438
rect 305102 706202 324546 706438
rect 324782 706202 324866 706438
rect 325102 706202 344546 706438
rect 344782 706202 344866 706438
rect 345102 706202 364546 706438
rect 364782 706202 364866 706438
rect 365102 706202 384546 706438
rect 384782 706202 384866 706438
rect 385102 706202 404546 706438
rect 404782 706202 404866 706438
rect 405102 706202 424546 706438
rect 424782 706202 424866 706438
rect 425102 706202 444546 706438
rect 444782 706202 444866 706438
rect 445102 706202 464546 706438
rect 464782 706202 464866 706438
rect 465102 706202 484546 706438
rect 484782 706202 484866 706438
rect 485102 706202 504546 706438
rect 504782 706202 504866 706438
rect 505102 706202 524546 706438
rect 524782 706202 524866 706438
rect 525102 706202 544546 706438
rect 544782 706202 544866 706438
rect 545102 706202 564546 706438
rect 564782 706202 564866 706438
rect 565102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 10826 705798
rect 11062 705562 11146 705798
rect 11382 705562 30826 705798
rect 31062 705562 31146 705798
rect 31382 705562 50826 705798
rect 51062 705562 51146 705798
rect 51382 705562 70826 705798
rect 71062 705562 71146 705798
rect 71382 705562 90826 705798
rect 91062 705562 91146 705798
rect 91382 705562 110826 705798
rect 111062 705562 111146 705798
rect 111382 705562 130826 705798
rect 131062 705562 131146 705798
rect 131382 705562 150826 705798
rect 151062 705562 151146 705798
rect 151382 705562 170826 705798
rect 171062 705562 171146 705798
rect 171382 705562 190826 705798
rect 191062 705562 191146 705798
rect 191382 705562 210826 705798
rect 211062 705562 211146 705798
rect 211382 705562 230826 705798
rect 231062 705562 231146 705798
rect 231382 705562 250826 705798
rect 251062 705562 251146 705798
rect 251382 705562 270826 705798
rect 271062 705562 271146 705798
rect 271382 705562 290826 705798
rect 291062 705562 291146 705798
rect 291382 705562 310826 705798
rect 311062 705562 311146 705798
rect 311382 705562 330826 705798
rect 331062 705562 331146 705798
rect 331382 705562 350826 705798
rect 351062 705562 351146 705798
rect 351382 705562 370826 705798
rect 371062 705562 371146 705798
rect 371382 705562 390826 705798
rect 391062 705562 391146 705798
rect 391382 705562 410826 705798
rect 411062 705562 411146 705798
rect 411382 705562 430826 705798
rect 431062 705562 431146 705798
rect 431382 705562 450826 705798
rect 451062 705562 451146 705798
rect 451382 705562 470826 705798
rect 471062 705562 471146 705798
rect 471382 705562 490826 705798
rect 491062 705562 491146 705798
rect 491382 705562 510826 705798
rect 511062 705562 511146 705798
rect 511382 705562 530826 705798
rect 531062 705562 531146 705798
rect 531382 705562 550826 705798
rect 551062 705562 551146 705798
rect 551382 705562 570826 705798
rect 571062 705562 571146 705798
rect 571382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 10826 705478
rect 11062 705242 11146 705478
rect 11382 705242 30826 705478
rect 31062 705242 31146 705478
rect 31382 705242 50826 705478
rect 51062 705242 51146 705478
rect 51382 705242 70826 705478
rect 71062 705242 71146 705478
rect 71382 705242 90826 705478
rect 91062 705242 91146 705478
rect 91382 705242 110826 705478
rect 111062 705242 111146 705478
rect 111382 705242 130826 705478
rect 131062 705242 131146 705478
rect 131382 705242 150826 705478
rect 151062 705242 151146 705478
rect 151382 705242 170826 705478
rect 171062 705242 171146 705478
rect 171382 705242 190826 705478
rect 191062 705242 191146 705478
rect 191382 705242 210826 705478
rect 211062 705242 211146 705478
rect 211382 705242 230826 705478
rect 231062 705242 231146 705478
rect 231382 705242 250826 705478
rect 251062 705242 251146 705478
rect 251382 705242 270826 705478
rect 271062 705242 271146 705478
rect 271382 705242 290826 705478
rect 291062 705242 291146 705478
rect 291382 705242 310826 705478
rect 311062 705242 311146 705478
rect 311382 705242 330826 705478
rect 331062 705242 331146 705478
rect 331382 705242 350826 705478
rect 351062 705242 351146 705478
rect 351382 705242 370826 705478
rect 371062 705242 371146 705478
rect 371382 705242 390826 705478
rect 391062 705242 391146 705478
rect 391382 705242 410826 705478
rect 411062 705242 411146 705478
rect 411382 705242 430826 705478
rect 431062 705242 431146 705478
rect 431382 705242 450826 705478
rect 451062 705242 451146 705478
rect 451382 705242 470826 705478
rect 471062 705242 471146 705478
rect 471382 705242 490826 705478
rect 491062 705242 491146 705478
rect 491382 705242 510826 705478
rect 511062 705242 511146 705478
rect 511382 705242 530826 705478
rect 531062 705242 531146 705478
rect 531382 705242 550826 705478
rect 551062 705242 551146 705478
rect 551382 705242 570826 705478
rect 571062 705242 571146 705478
rect 571382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 826 704838
rect 1062 704602 1146 704838
rect 1382 704602 20826 704838
rect 21062 704602 21146 704838
rect 21382 704602 40826 704838
rect 41062 704602 41146 704838
rect 41382 704602 60826 704838
rect 61062 704602 61146 704838
rect 61382 704602 80826 704838
rect 81062 704602 81146 704838
rect 81382 704602 100826 704838
rect 101062 704602 101146 704838
rect 101382 704602 120826 704838
rect 121062 704602 121146 704838
rect 121382 704602 140826 704838
rect 141062 704602 141146 704838
rect 141382 704602 160826 704838
rect 161062 704602 161146 704838
rect 161382 704602 180826 704838
rect 181062 704602 181146 704838
rect 181382 704602 200826 704838
rect 201062 704602 201146 704838
rect 201382 704602 220826 704838
rect 221062 704602 221146 704838
rect 221382 704602 240826 704838
rect 241062 704602 241146 704838
rect 241382 704602 260826 704838
rect 261062 704602 261146 704838
rect 261382 704602 280826 704838
rect 281062 704602 281146 704838
rect 281382 704602 300826 704838
rect 301062 704602 301146 704838
rect 301382 704602 320826 704838
rect 321062 704602 321146 704838
rect 321382 704602 340826 704838
rect 341062 704602 341146 704838
rect 341382 704602 360826 704838
rect 361062 704602 361146 704838
rect 361382 704602 380826 704838
rect 381062 704602 381146 704838
rect 381382 704602 400826 704838
rect 401062 704602 401146 704838
rect 401382 704602 420826 704838
rect 421062 704602 421146 704838
rect 421382 704602 440826 704838
rect 441062 704602 441146 704838
rect 441382 704602 460826 704838
rect 461062 704602 461146 704838
rect 461382 704602 480826 704838
rect 481062 704602 481146 704838
rect 481382 704602 500826 704838
rect 501062 704602 501146 704838
rect 501382 704602 520826 704838
rect 521062 704602 521146 704838
rect 521382 704602 540826 704838
rect 541062 704602 541146 704838
rect 541382 704602 560826 704838
rect 561062 704602 561146 704838
rect 561382 704602 580826 704838
rect 581062 704602 581146 704838
rect 581382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 826 704518
rect 1062 704282 1146 704518
rect 1382 704282 20826 704518
rect 21062 704282 21146 704518
rect 21382 704282 40826 704518
rect 41062 704282 41146 704518
rect 41382 704282 60826 704518
rect 61062 704282 61146 704518
rect 61382 704282 80826 704518
rect 81062 704282 81146 704518
rect 81382 704282 100826 704518
rect 101062 704282 101146 704518
rect 101382 704282 120826 704518
rect 121062 704282 121146 704518
rect 121382 704282 140826 704518
rect 141062 704282 141146 704518
rect 141382 704282 160826 704518
rect 161062 704282 161146 704518
rect 161382 704282 180826 704518
rect 181062 704282 181146 704518
rect 181382 704282 200826 704518
rect 201062 704282 201146 704518
rect 201382 704282 220826 704518
rect 221062 704282 221146 704518
rect 221382 704282 240826 704518
rect 241062 704282 241146 704518
rect 241382 704282 260826 704518
rect 261062 704282 261146 704518
rect 261382 704282 280826 704518
rect 281062 704282 281146 704518
rect 281382 704282 300826 704518
rect 301062 704282 301146 704518
rect 301382 704282 320826 704518
rect 321062 704282 321146 704518
rect 321382 704282 340826 704518
rect 341062 704282 341146 704518
rect 341382 704282 360826 704518
rect 361062 704282 361146 704518
rect 361382 704282 380826 704518
rect 381062 704282 381146 704518
rect 381382 704282 400826 704518
rect 401062 704282 401146 704518
rect 401382 704282 420826 704518
rect 421062 704282 421146 704518
rect 421382 704282 440826 704518
rect 441062 704282 441146 704518
rect 441382 704282 460826 704518
rect 461062 704282 461146 704518
rect 461382 704282 480826 704518
rect 481062 704282 481146 704518
rect 481382 704282 500826 704518
rect 501062 704282 501146 704518
rect 501382 704282 520826 704518
rect 521062 704282 521146 704518
rect 521382 704282 540826 704518
rect 541062 704282 541146 704518
rect 541382 704282 560826 704518
rect 561062 704282 561146 704518
rect 561382 704282 580826 704518
rect 581062 704282 581146 704518
rect 581382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 11986 698614
rect 12222 698378 12306 698614
rect 12542 698378 31986 698614
rect 32222 698378 32306 698614
rect 32542 698378 51986 698614
rect 52222 698378 52306 698614
rect 52542 698378 71986 698614
rect 72222 698378 72306 698614
rect 72542 698378 91986 698614
rect 92222 698378 92306 698614
rect 92542 698378 111986 698614
rect 112222 698378 112306 698614
rect 112542 698378 131986 698614
rect 132222 698378 132306 698614
rect 132542 698378 151986 698614
rect 152222 698378 152306 698614
rect 152542 698378 171986 698614
rect 172222 698378 172306 698614
rect 172542 698378 191986 698614
rect 192222 698378 192306 698614
rect 192542 698378 211986 698614
rect 212222 698378 212306 698614
rect 212542 698378 231986 698614
rect 232222 698378 232306 698614
rect 232542 698378 251986 698614
rect 252222 698378 252306 698614
rect 252542 698378 271986 698614
rect 272222 698378 272306 698614
rect 272542 698378 291986 698614
rect 292222 698378 292306 698614
rect 292542 698378 311986 698614
rect 312222 698378 312306 698614
rect 312542 698378 331986 698614
rect 332222 698378 332306 698614
rect 332542 698378 351986 698614
rect 352222 698378 352306 698614
rect 352542 698378 371986 698614
rect 372222 698378 372306 698614
rect 372542 698378 391986 698614
rect 392222 698378 392306 698614
rect 392542 698378 411986 698614
rect 412222 698378 412306 698614
rect 412542 698378 431986 698614
rect 432222 698378 432306 698614
rect 432542 698378 451986 698614
rect 452222 698378 452306 698614
rect 452542 698378 471986 698614
rect 472222 698378 472306 698614
rect 472542 698378 491986 698614
rect 492222 698378 492306 698614
rect 492542 698378 511986 698614
rect 512222 698378 512306 698614
rect 512542 698378 531986 698614
rect 532222 698378 532306 698614
rect 532542 698378 551986 698614
rect 552222 698378 552306 698614
rect 552542 698378 571986 698614
rect 572222 698378 572306 698614
rect 572542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 11986 698294
rect 12222 698058 12306 698294
rect 12542 698058 31986 698294
rect 32222 698058 32306 698294
rect 32542 698058 51986 698294
rect 52222 698058 52306 698294
rect 52542 698058 71986 698294
rect 72222 698058 72306 698294
rect 72542 698058 91986 698294
rect 92222 698058 92306 698294
rect 92542 698058 111986 698294
rect 112222 698058 112306 698294
rect 112542 698058 131986 698294
rect 132222 698058 132306 698294
rect 132542 698058 151986 698294
rect 152222 698058 152306 698294
rect 152542 698058 171986 698294
rect 172222 698058 172306 698294
rect 172542 698058 191986 698294
rect 192222 698058 192306 698294
rect 192542 698058 211986 698294
rect 212222 698058 212306 698294
rect 212542 698058 231986 698294
rect 232222 698058 232306 698294
rect 232542 698058 251986 698294
rect 252222 698058 252306 698294
rect 252542 698058 271986 698294
rect 272222 698058 272306 698294
rect 272542 698058 291986 698294
rect 292222 698058 292306 698294
rect 292542 698058 311986 698294
rect 312222 698058 312306 698294
rect 312542 698058 331986 698294
rect 332222 698058 332306 698294
rect 332542 698058 351986 698294
rect 352222 698058 352306 698294
rect 352542 698058 371986 698294
rect 372222 698058 372306 698294
rect 372542 698058 391986 698294
rect 392222 698058 392306 698294
rect 392542 698058 411986 698294
rect 412222 698058 412306 698294
rect 412542 698058 431986 698294
rect 432222 698058 432306 698294
rect 432542 698058 451986 698294
rect 452222 698058 452306 698294
rect 452542 698058 471986 698294
rect 472222 698058 472306 698294
rect 472542 698058 491986 698294
rect 492222 698058 492306 698294
rect 492542 698058 511986 698294
rect 512222 698058 512306 698294
rect 512542 698058 531986 698294
rect 532222 698058 532306 698294
rect 532542 698058 551986 698294
rect 552222 698058 552306 698294
rect 552542 698058 571986 698294
rect 572222 698058 572306 698294
rect 572542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 8266 694894
rect 8502 694658 8586 694894
rect 8822 694658 28266 694894
rect 28502 694658 28586 694894
rect 28822 694658 48266 694894
rect 48502 694658 48586 694894
rect 48822 694658 68266 694894
rect 68502 694658 68586 694894
rect 68822 694658 88266 694894
rect 88502 694658 88586 694894
rect 88822 694658 108266 694894
rect 108502 694658 108586 694894
rect 108822 694658 128266 694894
rect 128502 694658 128586 694894
rect 128822 694658 148266 694894
rect 148502 694658 148586 694894
rect 148822 694658 168266 694894
rect 168502 694658 168586 694894
rect 168822 694658 188266 694894
rect 188502 694658 188586 694894
rect 188822 694658 208266 694894
rect 208502 694658 208586 694894
rect 208822 694658 228266 694894
rect 228502 694658 228586 694894
rect 228822 694658 248266 694894
rect 248502 694658 248586 694894
rect 248822 694658 268266 694894
rect 268502 694658 268586 694894
rect 268822 694658 288266 694894
rect 288502 694658 288586 694894
rect 288822 694658 308266 694894
rect 308502 694658 308586 694894
rect 308822 694658 328266 694894
rect 328502 694658 328586 694894
rect 328822 694658 348266 694894
rect 348502 694658 348586 694894
rect 348822 694658 368266 694894
rect 368502 694658 368586 694894
rect 368822 694658 388266 694894
rect 388502 694658 388586 694894
rect 388822 694658 408266 694894
rect 408502 694658 408586 694894
rect 408822 694658 428266 694894
rect 428502 694658 428586 694894
rect 428822 694658 448266 694894
rect 448502 694658 448586 694894
rect 448822 694658 468266 694894
rect 468502 694658 468586 694894
rect 468822 694658 488266 694894
rect 488502 694658 488586 694894
rect 488822 694658 508266 694894
rect 508502 694658 508586 694894
rect 508822 694658 528266 694894
rect 528502 694658 528586 694894
rect 528822 694658 548266 694894
rect 548502 694658 548586 694894
rect 548822 694658 568266 694894
rect 568502 694658 568586 694894
rect 568822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 8266 694574
rect 8502 694338 8586 694574
rect 8822 694338 28266 694574
rect 28502 694338 28586 694574
rect 28822 694338 48266 694574
rect 48502 694338 48586 694574
rect 48822 694338 68266 694574
rect 68502 694338 68586 694574
rect 68822 694338 88266 694574
rect 88502 694338 88586 694574
rect 88822 694338 108266 694574
rect 108502 694338 108586 694574
rect 108822 694338 128266 694574
rect 128502 694338 128586 694574
rect 128822 694338 148266 694574
rect 148502 694338 148586 694574
rect 148822 694338 168266 694574
rect 168502 694338 168586 694574
rect 168822 694338 188266 694574
rect 188502 694338 188586 694574
rect 188822 694338 208266 694574
rect 208502 694338 208586 694574
rect 208822 694338 228266 694574
rect 228502 694338 228586 694574
rect 228822 694338 248266 694574
rect 248502 694338 248586 694574
rect 248822 694338 268266 694574
rect 268502 694338 268586 694574
rect 268822 694338 288266 694574
rect 288502 694338 288586 694574
rect 288822 694338 308266 694574
rect 308502 694338 308586 694574
rect 308822 694338 328266 694574
rect 328502 694338 328586 694574
rect 328822 694338 348266 694574
rect 348502 694338 348586 694574
rect 348822 694338 368266 694574
rect 368502 694338 368586 694574
rect 368822 694338 388266 694574
rect 388502 694338 388586 694574
rect 388822 694338 408266 694574
rect 408502 694338 408586 694574
rect 408822 694338 428266 694574
rect 428502 694338 428586 694574
rect 428822 694338 448266 694574
rect 448502 694338 448586 694574
rect 448822 694338 468266 694574
rect 468502 694338 468586 694574
rect 468822 694338 488266 694574
rect 488502 694338 488586 694574
rect 488822 694338 508266 694574
rect 508502 694338 508586 694574
rect 508822 694338 528266 694574
rect 528502 694338 528586 694574
rect 528822 694338 548266 694574
rect 548502 694338 548586 694574
rect 548822 694338 568266 694574
rect 568502 694338 568586 694574
rect 568822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 4546 691174
rect 4782 690938 4866 691174
rect 5102 690938 24546 691174
rect 24782 690938 24866 691174
rect 25102 690938 44546 691174
rect 44782 690938 44866 691174
rect 45102 690938 64546 691174
rect 64782 690938 64866 691174
rect 65102 690938 84546 691174
rect 84782 690938 84866 691174
rect 85102 690938 104546 691174
rect 104782 690938 104866 691174
rect 105102 690938 124546 691174
rect 124782 690938 124866 691174
rect 125102 690938 144546 691174
rect 144782 690938 144866 691174
rect 145102 690938 164546 691174
rect 164782 690938 164866 691174
rect 165102 690938 184546 691174
rect 184782 690938 184866 691174
rect 185102 690938 204546 691174
rect 204782 690938 204866 691174
rect 205102 690938 224546 691174
rect 224782 690938 224866 691174
rect 225102 690938 244546 691174
rect 244782 690938 244866 691174
rect 245102 690938 264546 691174
rect 264782 690938 264866 691174
rect 265102 690938 284546 691174
rect 284782 690938 284866 691174
rect 285102 690938 304546 691174
rect 304782 690938 304866 691174
rect 305102 690938 324546 691174
rect 324782 690938 324866 691174
rect 325102 690938 344546 691174
rect 344782 690938 344866 691174
rect 345102 690938 364546 691174
rect 364782 690938 364866 691174
rect 365102 690938 384546 691174
rect 384782 690938 384866 691174
rect 385102 690938 404546 691174
rect 404782 690938 404866 691174
rect 405102 690938 424546 691174
rect 424782 690938 424866 691174
rect 425102 690938 444546 691174
rect 444782 690938 444866 691174
rect 445102 690938 464546 691174
rect 464782 690938 464866 691174
rect 465102 690938 484546 691174
rect 484782 690938 484866 691174
rect 485102 690938 504546 691174
rect 504782 690938 504866 691174
rect 505102 690938 524546 691174
rect 524782 690938 524866 691174
rect 525102 690938 544546 691174
rect 544782 690938 544866 691174
rect 545102 690938 564546 691174
rect 564782 690938 564866 691174
rect 565102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 4546 690854
rect 4782 690618 4866 690854
rect 5102 690618 24546 690854
rect 24782 690618 24866 690854
rect 25102 690618 44546 690854
rect 44782 690618 44866 690854
rect 45102 690618 64546 690854
rect 64782 690618 64866 690854
rect 65102 690618 84546 690854
rect 84782 690618 84866 690854
rect 85102 690618 104546 690854
rect 104782 690618 104866 690854
rect 105102 690618 124546 690854
rect 124782 690618 124866 690854
rect 125102 690618 144546 690854
rect 144782 690618 144866 690854
rect 145102 690618 164546 690854
rect 164782 690618 164866 690854
rect 165102 690618 184546 690854
rect 184782 690618 184866 690854
rect 185102 690618 204546 690854
rect 204782 690618 204866 690854
rect 205102 690618 224546 690854
rect 224782 690618 224866 690854
rect 225102 690618 244546 690854
rect 244782 690618 244866 690854
rect 245102 690618 264546 690854
rect 264782 690618 264866 690854
rect 265102 690618 284546 690854
rect 284782 690618 284866 690854
rect 285102 690618 304546 690854
rect 304782 690618 304866 690854
rect 305102 690618 324546 690854
rect 324782 690618 324866 690854
rect 325102 690618 344546 690854
rect 344782 690618 344866 690854
rect 345102 690618 364546 690854
rect 364782 690618 364866 690854
rect 365102 690618 384546 690854
rect 384782 690618 384866 690854
rect 385102 690618 404546 690854
rect 404782 690618 404866 690854
rect 405102 690618 424546 690854
rect 424782 690618 424866 690854
rect 425102 690618 444546 690854
rect 444782 690618 444866 690854
rect 445102 690618 464546 690854
rect 464782 690618 464866 690854
rect 465102 690618 484546 690854
rect 484782 690618 484866 690854
rect 485102 690618 504546 690854
rect 504782 690618 504866 690854
rect 505102 690618 524546 690854
rect 524782 690618 524866 690854
rect 525102 690618 544546 690854
rect 544782 690618 544866 690854
rect 545102 690618 564546 690854
rect 564782 690618 564866 690854
rect 565102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 826 687454
rect 1062 687218 1146 687454
rect 1382 687218 20826 687454
rect 21062 687218 21146 687454
rect 21382 687218 40826 687454
rect 41062 687218 41146 687454
rect 41382 687218 60826 687454
rect 61062 687218 61146 687454
rect 61382 687218 80826 687454
rect 81062 687218 81146 687454
rect 81382 687218 100826 687454
rect 101062 687218 101146 687454
rect 101382 687218 120826 687454
rect 121062 687218 121146 687454
rect 121382 687218 140826 687454
rect 141062 687218 141146 687454
rect 141382 687218 160826 687454
rect 161062 687218 161146 687454
rect 161382 687218 180826 687454
rect 181062 687218 181146 687454
rect 181382 687218 200826 687454
rect 201062 687218 201146 687454
rect 201382 687218 220826 687454
rect 221062 687218 221146 687454
rect 221382 687218 240826 687454
rect 241062 687218 241146 687454
rect 241382 687218 260826 687454
rect 261062 687218 261146 687454
rect 261382 687218 280826 687454
rect 281062 687218 281146 687454
rect 281382 687218 300826 687454
rect 301062 687218 301146 687454
rect 301382 687218 320826 687454
rect 321062 687218 321146 687454
rect 321382 687218 340826 687454
rect 341062 687218 341146 687454
rect 341382 687218 360826 687454
rect 361062 687218 361146 687454
rect 361382 687218 380826 687454
rect 381062 687218 381146 687454
rect 381382 687218 400826 687454
rect 401062 687218 401146 687454
rect 401382 687218 420826 687454
rect 421062 687218 421146 687454
rect 421382 687218 440826 687454
rect 441062 687218 441146 687454
rect 441382 687218 460826 687454
rect 461062 687218 461146 687454
rect 461382 687218 480826 687454
rect 481062 687218 481146 687454
rect 481382 687218 500826 687454
rect 501062 687218 501146 687454
rect 501382 687218 520826 687454
rect 521062 687218 521146 687454
rect 521382 687218 540826 687454
rect 541062 687218 541146 687454
rect 541382 687218 560826 687454
rect 561062 687218 561146 687454
rect 561382 687218 580826 687454
rect 581062 687218 581146 687454
rect 581382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 826 687134
rect 1062 686898 1146 687134
rect 1382 686898 20826 687134
rect 21062 686898 21146 687134
rect 21382 686898 40826 687134
rect 41062 686898 41146 687134
rect 41382 686898 60826 687134
rect 61062 686898 61146 687134
rect 61382 686898 80826 687134
rect 81062 686898 81146 687134
rect 81382 686898 100826 687134
rect 101062 686898 101146 687134
rect 101382 686898 120826 687134
rect 121062 686898 121146 687134
rect 121382 686898 140826 687134
rect 141062 686898 141146 687134
rect 141382 686898 160826 687134
rect 161062 686898 161146 687134
rect 161382 686898 180826 687134
rect 181062 686898 181146 687134
rect 181382 686898 200826 687134
rect 201062 686898 201146 687134
rect 201382 686898 220826 687134
rect 221062 686898 221146 687134
rect 221382 686898 240826 687134
rect 241062 686898 241146 687134
rect 241382 686898 260826 687134
rect 261062 686898 261146 687134
rect 261382 686898 280826 687134
rect 281062 686898 281146 687134
rect 281382 686898 300826 687134
rect 301062 686898 301146 687134
rect 301382 686898 320826 687134
rect 321062 686898 321146 687134
rect 321382 686898 340826 687134
rect 341062 686898 341146 687134
rect 341382 686898 360826 687134
rect 361062 686898 361146 687134
rect 361382 686898 380826 687134
rect 381062 686898 381146 687134
rect 381382 686898 400826 687134
rect 401062 686898 401146 687134
rect 401382 686898 420826 687134
rect 421062 686898 421146 687134
rect 421382 686898 440826 687134
rect 441062 686898 441146 687134
rect 441382 686898 460826 687134
rect 461062 686898 461146 687134
rect 461382 686898 480826 687134
rect 481062 686898 481146 687134
rect 481382 686898 500826 687134
rect 501062 686898 501146 687134
rect 501382 686898 520826 687134
rect 521062 686898 521146 687134
rect 521382 686898 540826 687134
rect 541062 686898 541146 687134
rect 541382 686898 560826 687134
rect 561062 686898 561146 687134
rect 561382 686898 580826 687134
rect 581062 686898 581146 687134
rect 581382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 21986 680614
rect 22222 680378 22306 680614
rect 22542 680378 41986 680614
rect 42222 680378 42306 680614
rect 42542 680378 61986 680614
rect 62222 680378 62306 680614
rect 62542 680378 81986 680614
rect 82222 680378 82306 680614
rect 82542 680378 101986 680614
rect 102222 680378 102306 680614
rect 102542 680378 121986 680614
rect 122222 680378 122306 680614
rect 122542 680378 141986 680614
rect 142222 680378 142306 680614
rect 142542 680378 161986 680614
rect 162222 680378 162306 680614
rect 162542 680378 181986 680614
rect 182222 680378 182306 680614
rect 182542 680378 201986 680614
rect 202222 680378 202306 680614
rect 202542 680378 221986 680614
rect 222222 680378 222306 680614
rect 222542 680378 241986 680614
rect 242222 680378 242306 680614
rect 242542 680378 261986 680614
rect 262222 680378 262306 680614
rect 262542 680378 281986 680614
rect 282222 680378 282306 680614
rect 282542 680378 301986 680614
rect 302222 680378 302306 680614
rect 302542 680378 321986 680614
rect 322222 680378 322306 680614
rect 322542 680378 341986 680614
rect 342222 680378 342306 680614
rect 342542 680378 361986 680614
rect 362222 680378 362306 680614
rect 362542 680378 381986 680614
rect 382222 680378 382306 680614
rect 382542 680378 401986 680614
rect 402222 680378 402306 680614
rect 402542 680378 421986 680614
rect 422222 680378 422306 680614
rect 422542 680378 441986 680614
rect 442222 680378 442306 680614
rect 442542 680378 461986 680614
rect 462222 680378 462306 680614
rect 462542 680378 481986 680614
rect 482222 680378 482306 680614
rect 482542 680378 501986 680614
rect 502222 680378 502306 680614
rect 502542 680378 521986 680614
rect 522222 680378 522306 680614
rect 522542 680378 541986 680614
rect 542222 680378 542306 680614
rect 542542 680378 561986 680614
rect 562222 680378 562306 680614
rect 562542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 21986 680294
rect 22222 680058 22306 680294
rect 22542 680058 41986 680294
rect 42222 680058 42306 680294
rect 42542 680058 61986 680294
rect 62222 680058 62306 680294
rect 62542 680058 81986 680294
rect 82222 680058 82306 680294
rect 82542 680058 101986 680294
rect 102222 680058 102306 680294
rect 102542 680058 121986 680294
rect 122222 680058 122306 680294
rect 122542 680058 141986 680294
rect 142222 680058 142306 680294
rect 142542 680058 161986 680294
rect 162222 680058 162306 680294
rect 162542 680058 181986 680294
rect 182222 680058 182306 680294
rect 182542 680058 201986 680294
rect 202222 680058 202306 680294
rect 202542 680058 221986 680294
rect 222222 680058 222306 680294
rect 222542 680058 241986 680294
rect 242222 680058 242306 680294
rect 242542 680058 261986 680294
rect 262222 680058 262306 680294
rect 262542 680058 281986 680294
rect 282222 680058 282306 680294
rect 282542 680058 301986 680294
rect 302222 680058 302306 680294
rect 302542 680058 321986 680294
rect 322222 680058 322306 680294
rect 322542 680058 341986 680294
rect 342222 680058 342306 680294
rect 342542 680058 361986 680294
rect 362222 680058 362306 680294
rect 362542 680058 381986 680294
rect 382222 680058 382306 680294
rect 382542 680058 401986 680294
rect 402222 680058 402306 680294
rect 402542 680058 421986 680294
rect 422222 680058 422306 680294
rect 422542 680058 441986 680294
rect 442222 680058 442306 680294
rect 442542 680058 461986 680294
rect 462222 680058 462306 680294
rect 462542 680058 481986 680294
rect 482222 680058 482306 680294
rect 482542 680058 501986 680294
rect 502222 680058 502306 680294
rect 502542 680058 521986 680294
rect 522222 680058 522306 680294
rect 522542 680058 541986 680294
rect 542222 680058 542306 680294
rect 542542 680058 561986 680294
rect 562222 680058 562306 680294
rect 562542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 18266 676894
rect 18502 676658 18586 676894
rect 18822 676658 38266 676894
rect 38502 676658 38586 676894
rect 38822 676658 58266 676894
rect 58502 676658 58586 676894
rect 58822 676658 78266 676894
rect 78502 676658 78586 676894
rect 78822 676658 98266 676894
rect 98502 676658 98586 676894
rect 98822 676658 118266 676894
rect 118502 676658 118586 676894
rect 118822 676658 138266 676894
rect 138502 676658 138586 676894
rect 138822 676658 158266 676894
rect 158502 676658 158586 676894
rect 158822 676658 178266 676894
rect 178502 676658 178586 676894
rect 178822 676658 198266 676894
rect 198502 676658 198586 676894
rect 198822 676658 218266 676894
rect 218502 676658 218586 676894
rect 218822 676658 238266 676894
rect 238502 676658 238586 676894
rect 238822 676658 258266 676894
rect 258502 676658 258586 676894
rect 258822 676658 278266 676894
rect 278502 676658 278586 676894
rect 278822 676658 298266 676894
rect 298502 676658 298586 676894
rect 298822 676658 318266 676894
rect 318502 676658 318586 676894
rect 318822 676658 338266 676894
rect 338502 676658 338586 676894
rect 338822 676658 358266 676894
rect 358502 676658 358586 676894
rect 358822 676658 378266 676894
rect 378502 676658 378586 676894
rect 378822 676658 398266 676894
rect 398502 676658 398586 676894
rect 398822 676658 418266 676894
rect 418502 676658 418586 676894
rect 418822 676658 438266 676894
rect 438502 676658 438586 676894
rect 438822 676658 458266 676894
rect 458502 676658 458586 676894
rect 458822 676658 478266 676894
rect 478502 676658 478586 676894
rect 478822 676658 498266 676894
rect 498502 676658 498586 676894
rect 498822 676658 518266 676894
rect 518502 676658 518586 676894
rect 518822 676658 538266 676894
rect 538502 676658 538586 676894
rect 538822 676658 558266 676894
rect 558502 676658 558586 676894
rect 558822 676658 578266 676894
rect 578502 676658 578586 676894
rect 578822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 18266 676574
rect 18502 676338 18586 676574
rect 18822 676338 38266 676574
rect 38502 676338 38586 676574
rect 38822 676338 58266 676574
rect 58502 676338 58586 676574
rect 58822 676338 78266 676574
rect 78502 676338 78586 676574
rect 78822 676338 98266 676574
rect 98502 676338 98586 676574
rect 98822 676338 118266 676574
rect 118502 676338 118586 676574
rect 118822 676338 138266 676574
rect 138502 676338 138586 676574
rect 138822 676338 158266 676574
rect 158502 676338 158586 676574
rect 158822 676338 178266 676574
rect 178502 676338 178586 676574
rect 178822 676338 198266 676574
rect 198502 676338 198586 676574
rect 198822 676338 218266 676574
rect 218502 676338 218586 676574
rect 218822 676338 238266 676574
rect 238502 676338 238586 676574
rect 238822 676338 258266 676574
rect 258502 676338 258586 676574
rect 258822 676338 278266 676574
rect 278502 676338 278586 676574
rect 278822 676338 298266 676574
rect 298502 676338 298586 676574
rect 298822 676338 318266 676574
rect 318502 676338 318586 676574
rect 318822 676338 338266 676574
rect 338502 676338 338586 676574
rect 338822 676338 358266 676574
rect 358502 676338 358586 676574
rect 358822 676338 378266 676574
rect 378502 676338 378586 676574
rect 378822 676338 398266 676574
rect 398502 676338 398586 676574
rect 398822 676338 418266 676574
rect 418502 676338 418586 676574
rect 418822 676338 438266 676574
rect 438502 676338 438586 676574
rect 438822 676338 458266 676574
rect 458502 676338 458586 676574
rect 458822 676338 478266 676574
rect 478502 676338 478586 676574
rect 478822 676338 498266 676574
rect 498502 676338 498586 676574
rect 498822 676338 518266 676574
rect 518502 676338 518586 676574
rect 518822 676338 538266 676574
rect 538502 676338 538586 676574
rect 538822 676338 558266 676574
rect 558502 676338 558586 676574
rect 558822 676338 578266 676574
rect 578502 676338 578586 676574
rect 578822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 14546 673174
rect 14782 672938 14866 673174
rect 15102 672938 34546 673174
rect 34782 672938 34866 673174
rect 35102 672938 54546 673174
rect 54782 672938 54866 673174
rect 55102 672938 74546 673174
rect 74782 672938 74866 673174
rect 75102 672938 94546 673174
rect 94782 672938 94866 673174
rect 95102 672938 114546 673174
rect 114782 672938 114866 673174
rect 115102 672938 134546 673174
rect 134782 672938 134866 673174
rect 135102 672938 154546 673174
rect 154782 672938 154866 673174
rect 155102 672938 174546 673174
rect 174782 672938 174866 673174
rect 175102 672938 194546 673174
rect 194782 672938 194866 673174
rect 195102 672938 214546 673174
rect 214782 672938 214866 673174
rect 215102 672938 234546 673174
rect 234782 672938 234866 673174
rect 235102 672938 254546 673174
rect 254782 672938 254866 673174
rect 255102 672938 274546 673174
rect 274782 672938 274866 673174
rect 275102 672938 294546 673174
rect 294782 672938 294866 673174
rect 295102 672938 314546 673174
rect 314782 672938 314866 673174
rect 315102 672938 334546 673174
rect 334782 672938 334866 673174
rect 335102 672938 354546 673174
rect 354782 672938 354866 673174
rect 355102 672938 374546 673174
rect 374782 672938 374866 673174
rect 375102 672938 394546 673174
rect 394782 672938 394866 673174
rect 395102 672938 414546 673174
rect 414782 672938 414866 673174
rect 415102 672938 434546 673174
rect 434782 672938 434866 673174
rect 435102 672938 454546 673174
rect 454782 672938 454866 673174
rect 455102 672938 474546 673174
rect 474782 672938 474866 673174
rect 475102 672938 494546 673174
rect 494782 672938 494866 673174
rect 495102 672938 514546 673174
rect 514782 672938 514866 673174
rect 515102 672938 534546 673174
rect 534782 672938 534866 673174
rect 535102 672938 554546 673174
rect 554782 672938 554866 673174
rect 555102 672938 574546 673174
rect 574782 672938 574866 673174
rect 575102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 14546 672854
rect 14782 672618 14866 672854
rect 15102 672618 34546 672854
rect 34782 672618 34866 672854
rect 35102 672618 54546 672854
rect 54782 672618 54866 672854
rect 55102 672618 74546 672854
rect 74782 672618 74866 672854
rect 75102 672618 94546 672854
rect 94782 672618 94866 672854
rect 95102 672618 114546 672854
rect 114782 672618 114866 672854
rect 115102 672618 134546 672854
rect 134782 672618 134866 672854
rect 135102 672618 154546 672854
rect 154782 672618 154866 672854
rect 155102 672618 174546 672854
rect 174782 672618 174866 672854
rect 175102 672618 194546 672854
rect 194782 672618 194866 672854
rect 195102 672618 214546 672854
rect 214782 672618 214866 672854
rect 215102 672618 234546 672854
rect 234782 672618 234866 672854
rect 235102 672618 254546 672854
rect 254782 672618 254866 672854
rect 255102 672618 274546 672854
rect 274782 672618 274866 672854
rect 275102 672618 294546 672854
rect 294782 672618 294866 672854
rect 295102 672618 314546 672854
rect 314782 672618 314866 672854
rect 315102 672618 334546 672854
rect 334782 672618 334866 672854
rect 335102 672618 354546 672854
rect 354782 672618 354866 672854
rect 355102 672618 374546 672854
rect 374782 672618 374866 672854
rect 375102 672618 394546 672854
rect 394782 672618 394866 672854
rect 395102 672618 414546 672854
rect 414782 672618 414866 672854
rect 415102 672618 434546 672854
rect 434782 672618 434866 672854
rect 435102 672618 454546 672854
rect 454782 672618 454866 672854
rect 455102 672618 474546 672854
rect 474782 672618 474866 672854
rect 475102 672618 494546 672854
rect 494782 672618 494866 672854
rect 495102 672618 514546 672854
rect 514782 672618 514866 672854
rect 515102 672618 534546 672854
rect 534782 672618 534866 672854
rect 535102 672618 554546 672854
rect 554782 672618 554866 672854
rect 555102 672618 574546 672854
rect 574782 672618 574866 672854
rect 575102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 10826 669454
rect 11062 669218 11146 669454
rect 11382 669218 30826 669454
rect 31062 669218 31146 669454
rect 31382 669218 50826 669454
rect 51062 669218 51146 669454
rect 51382 669218 70826 669454
rect 71062 669218 71146 669454
rect 71382 669218 90826 669454
rect 91062 669218 91146 669454
rect 91382 669218 110826 669454
rect 111062 669218 111146 669454
rect 111382 669218 130826 669454
rect 131062 669218 131146 669454
rect 131382 669218 150826 669454
rect 151062 669218 151146 669454
rect 151382 669218 170826 669454
rect 171062 669218 171146 669454
rect 171382 669218 190826 669454
rect 191062 669218 191146 669454
rect 191382 669218 210826 669454
rect 211062 669218 211146 669454
rect 211382 669218 230826 669454
rect 231062 669218 231146 669454
rect 231382 669218 250826 669454
rect 251062 669218 251146 669454
rect 251382 669218 270826 669454
rect 271062 669218 271146 669454
rect 271382 669218 290826 669454
rect 291062 669218 291146 669454
rect 291382 669218 310826 669454
rect 311062 669218 311146 669454
rect 311382 669218 330826 669454
rect 331062 669218 331146 669454
rect 331382 669218 350826 669454
rect 351062 669218 351146 669454
rect 351382 669218 370826 669454
rect 371062 669218 371146 669454
rect 371382 669218 390826 669454
rect 391062 669218 391146 669454
rect 391382 669218 410826 669454
rect 411062 669218 411146 669454
rect 411382 669218 430826 669454
rect 431062 669218 431146 669454
rect 431382 669218 450826 669454
rect 451062 669218 451146 669454
rect 451382 669218 470826 669454
rect 471062 669218 471146 669454
rect 471382 669218 490826 669454
rect 491062 669218 491146 669454
rect 491382 669218 510826 669454
rect 511062 669218 511146 669454
rect 511382 669218 530826 669454
rect 531062 669218 531146 669454
rect 531382 669218 550826 669454
rect 551062 669218 551146 669454
rect 551382 669218 570826 669454
rect 571062 669218 571146 669454
rect 571382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 10826 669134
rect 11062 668898 11146 669134
rect 11382 668898 30826 669134
rect 31062 668898 31146 669134
rect 31382 668898 50826 669134
rect 51062 668898 51146 669134
rect 51382 668898 70826 669134
rect 71062 668898 71146 669134
rect 71382 668898 90826 669134
rect 91062 668898 91146 669134
rect 91382 668898 110826 669134
rect 111062 668898 111146 669134
rect 111382 668898 130826 669134
rect 131062 668898 131146 669134
rect 131382 668898 150826 669134
rect 151062 668898 151146 669134
rect 151382 668898 170826 669134
rect 171062 668898 171146 669134
rect 171382 668898 190826 669134
rect 191062 668898 191146 669134
rect 191382 668898 210826 669134
rect 211062 668898 211146 669134
rect 211382 668898 230826 669134
rect 231062 668898 231146 669134
rect 231382 668898 250826 669134
rect 251062 668898 251146 669134
rect 251382 668898 270826 669134
rect 271062 668898 271146 669134
rect 271382 668898 290826 669134
rect 291062 668898 291146 669134
rect 291382 668898 310826 669134
rect 311062 668898 311146 669134
rect 311382 668898 330826 669134
rect 331062 668898 331146 669134
rect 331382 668898 350826 669134
rect 351062 668898 351146 669134
rect 351382 668898 370826 669134
rect 371062 668898 371146 669134
rect 371382 668898 390826 669134
rect 391062 668898 391146 669134
rect 391382 668898 410826 669134
rect 411062 668898 411146 669134
rect 411382 668898 430826 669134
rect 431062 668898 431146 669134
rect 431382 668898 450826 669134
rect 451062 668898 451146 669134
rect 451382 668898 470826 669134
rect 471062 668898 471146 669134
rect 471382 668898 490826 669134
rect 491062 668898 491146 669134
rect 491382 668898 510826 669134
rect 511062 668898 511146 669134
rect 511382 668898 530826 669134
rect 531062 668898 531146 669134
rect 531382 668898 550826 669134
rect 551062 668898 551146 669134
rect 551382 668898 570826 669134
rect 571062 668898 571146 669134
rect 571382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 11986 662614
rect 12222 662378 12306 662614
rect 12542 662378 31986 662614
rect 32222 662378 32306 662614
rect 32542 662378 51986 662614
rect 52222 662378 52306 662614
rect 52542 662378 71986 662614
rect 72222 662378 72306 662614
rect 72542 662378 91986 662614
rect 92222 662378 92306 662614
rect 92542 662378 111986 662614
rect 112222 662378 112306 662614
rect 112542 662378 131986 662614
rect 132222 662378 132306 662614
rect 132542 662378 151986 662614
rect 152222 662378 152306 662614
rect 152542 662378 171986 662614
rect 172222 662378 172306 662614
rect 172542 662378 191986 662614
rect 192222 662378 192306 662614
rect 192542 662378 211986 662614
rect 212222 662378 212306 662614
rect 212542 662378 231986 662614
rect 232222 662378 232306 662614
rect 232542 662378 251986 662614
rect 252222 662378 252306 662614
rect 252542 662378 271986 662614
rect 272222 662378 272306 662614
rect 272542 662378 291986 662614
rect 292222 662378 292306 662614
rect 292542 662378 311986 662614
rect 312222 662378 312306 662614
rect 312542 662378 331986 662614
rect 332222 662378 332306 662614
rect 332542 662378 351986 662614
rect 352222 662378 352306 662614
rect 352542 662378 371986 662614
rect 372222 662378 372306 662614
rect 372542 662378 391986 662614
rect 392222 662378 392306 662614
rect 392542 662378 411986 662614
rect 412222 662378 412306 662614
rect 412542 662378 431986 662614
rect 432222 662378 432306 662614
rect 432542 662378 451986 662614
rect 452222 662378 452306 662614
rect 452542 662378 471986 662614
rect 472222 662378 472306 662614
rect 472542 662378 491986 662614
rect 492222 662378 492306 662614
rect 492542 662378 511986 662614
rect 512222 662378 512306 662614
rect 512542 662378 531986 662614
rect 532222 662378 532306 662614
rect 532542 662378 551986 662614
rect 552222 662378 552306 662614
rect 552542 662378 571986 662614
rect 572222 662378 572306 662614
rect 572542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 11986 662294
rect 12222 662058 12306 662294
rect 12542 662058 31986 662294
rect 32222 662058 32306 662294
rect 32542 662058 51986 662294
rect 52222 662058 52306 662294
rect 52542 662058 71986 662294
rect 72222 662058 72306 662294
rect 72542 662058 91986 662294
rect 92222 662058 92306 662294
rect 92542 662058 111986 662294
rect 112222 662058 112306 662294
rect 112542 662058 131986 662294
rect 132222 662058 132306 662294
rect 132542 662058 151986 662294
rect 152222 662058 152306 662294
rect 152542 662058 171986 662294
rect 172222 662058 172306 662294
rect 172542 662058 191986 662294
rect 192222 662058 192306 662294
rect 192542 662058 211986 662294
rect 212222 662058 212306 662294
rect 212542 662058 231986 662294
rect 232222 662058 232306 662294
rect 232542 662058 251986 662294
rect 252222 662058 252306 662294
rect 252542 662058 271986 662294
rect 272222 662058 272306 662294
rect 272542 662058 291986 662294
rect 292222 662058 292306 662294
rect 292542 662058 311986 662294
rect 312222 662058 312306 662294
rect 312542 662058 331986 662294
rect 332222 662058 332306 662294
rect 332542 662058 351986 662294
rect 352222 662058 352306 662294
rect 352542 662058 371986 662294
rect 372222 662058 372306 662294
rect 372542 662058 391986 662294
rect 392222 662058 392306 662294
rect 392542 662058 411986 662294
rect 412222 662058 412306 662294
rect 412542 662058 431986 662294
rect 432222 662058 432306 662294
rect 432542 662058 451986 662294
rect 452222 662058 452306 662294
rect 452542 662058 471986 662294
rect 472222 662058 472306 662294
rect 472542 662058 491986 662294
rect 492222 662058 492306 662294
rect 492542 662058 511986 662294
rect 512222 662058 512306 662294
rect 512542 662058 531986 662294
rect 532222 662058 532306 662294
rect 532542 662058 551986 662294
rect 552222 662058 552306 662294
rect 552542 662058 571986 662294
rect 572222 662058 572306 662294
rect 572542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 8266 658894
rect 8502 658658 8586 658894
rect 8822 658658 28266 658894
rect 28502 658658 28586 658894
rect 28822 658658 48266 658894
rect 48502 658658 48586 658894
rect 48822 658658 68266 658894
rect 68502 658658 68586 658894
rect 68822 658658 88266 658894
rect 88502 658658 88586 658894
rect 88822 658658 108266 658894
rect 108502 658658 108586 658894
rect 108822 658658 128266 658894
rect 128502 658658 128586 658894
rect 128822 658658 148266 658894
rect 148502 658658 148586 658894
rect 148822 658658 168266 658894
rect 168502 658658 168586 658894
rect 168822 658658 188266 658894
rect 188502 658658 188586 658894
rect 188822 658658 208266 658894
rect 208502 658658 208586 658894
rect 208822 658658 228266 658894
rect 228502 658658 228586 658894
rect 228822 658658 248266 658894
rect 248502 658658 248586 658894
rect 248822 658658 268266 658894
rect 268502 658658 268586 658894
rect 268822 658658 288266 658894
rect 288502 658658 288586 658894
rect 288822 658658 308266 658894
rect 308502 658658 308586 658894
rect 308822 658658 328266 658894
rect 328502 658658 328586 658894
rect 328822 658658 348266 658894
rect 348502 658658 348586 658894
rect 348822 658658 368266 658894
rect 368502 658658 368586 658894
rect 368822 658658 388266 658894
rect 388502 658658 388586 658894
rect 388822 658658 408266 658894
rect 408502 658658 408586 658894
rect 408822 658658 428266 658894
rect 428502 658658 428586 658894
rect 428822 658658 448266 658894
rect 448502 658658 448586 658894
rect 448822 658658 468266 658894
rect 468502 658658 468586 658894
rect 468822 658658 488266 658894
rect 488502 658658 488586 658894
rect 488822 658658 508266 658894
rect 508502 658658 508586 658894
rect 508822 658658 528266 658894
rect 528502 658658 528586 658894
rect 528822 658658 548266 658894
rect 548502 658658 548586 658894
rect 548822 658658 568266 658894
rect 568502 658658 568586 658894
rect 568822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 8266 658574
rect 8502 658338 8586 658574
rect 8822 658338 28266 658574
rect 28502 658338 28586 658574
rect 28822 658338 48266 658574
rect 48502 658338 48586 658574
rect 48822 658338 68266 658574
rect 68502 658338 68586 658574
rect 68822 658338 88266 658574
rect 88502 658338 88586 658574
rect 88822 658338 108266 658574
rect 108502 658338 108586 658574
rect 108822 658338 128266 658574
rect 128502 658338 128586 658574
rect 128822 658338 148266 658574
rect 148502 658338 148586 658574
rect 148822 658338 168266 658574
rect 168502 658338 168586 658574
rect 168822 658338 188266 658574
rect 188502 658338 188586 658574
rect 188822 658338 208266 658574
rect 208502 658338 208586 658574
rect 208822 658338 228266 658574
rect 228502 658338 228586 658574
rect 228822 658338 248266 658574
rect 248502 658338 248586 658574
rect 248822 658338 268266 658574
rect 268502 658338 268586 658574
rect 268822 658338 288266 658574
rect 288502 658338 288586 658574
rect 288822 658338 308266 658574
rect 308502 658338 308586 658574
rect 308822 658338 328266 658574
rect 328502 658338 328586 658574
rect 328822 658338 348266 658574
rect 348502 658338 348586 658574
rect 348822 658338 368266 658574
rect 368502 658338 368586 658574
rect 368822 658338 388266 658574
rect 388502 658338 388586 658574
rect 388822 658338 408266 658574
rect 408502 658338 408586 658574
rect 408822 658338 428266 658574
rect 428502 658338 428586 658574
rect 428822 658338 448266 658574
rect 448502 658338 448586 658574
rect 448822 658338 468266 658574
rect 468502 658338 468586 658574
rect 468822 658338 488266 658574
rect 488502 658338 488586 658574
rect 488822 658338 508266 658574
rect 508502 658338 508586 658574
rect 508822 658338 528266 658574
rect 528502 658338 528586 658574
rect 528822 658338 548266 658574
rect 548502 658338 548586 658574
rect 548822 658338 568266 658574
rect 568502 658338 568586 658574
rect 568822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 4546 655174
rect 4782 654938 4866 655174
rect 5102 654938 24546 655174
rect 24782 654938 24866 655174
rect 25102 654938 44546 655174
rect 44782 654938 44866 655174
rect 45102 654938 64546 655174
rect 64782 654938 64866 655174
rect 65102 654938 84546 655174
rect 84782 654938 84866 655174
rect 85102 654938 104546 655174
rect 104782 654938 104866 655174
rect 105102 654938 124546 655174
rect 124782 654938 124866 655174
rect 125102 654938 144546 655174
rect 144782 654938 144866 655174
rect 145102 654938 164546 655174
rect 164782 654938 164866 655174
rect 165102 654938 184546 655174
rect 184782 654938 184866 655174
rect 185102 654938 204546 655174
rect 204782 654938 204866 655174
rect 205102 654938 224546 655174
rect 224782 654938 224866 655174
rect 225102 654938 244546 655174
rect 244782 654938 244866 655174
rect 245102 654938 264546 655174
rect 264782 654938 264866 655174
rect 265102 654938 284546 655174
rect 284782 654938 284866 655174
rect 285102 654938 304546 655174
rect 304782 654938 304866 655174
rect 305102 654938 324546 655174
rect 324782 654938 324866 655174
rect 325102 654938 344546 655174
rect 344782 654938 344866 655174
rect 345102 654938 364546 655174
rect 364782 654938 364866 655174
rect 365102 654938 384546 655174
rect 384782 654938 384866 655174
rect 385102 654938 404546 655174
rect 404782 654938 404866 655174
rect 405102 654938 424546 655174
rect 424782 654938 424866 655174
rect 425102 654938 444546 655174
rect 444782 654938 444866 655174
rect 445102 654938 464546 655174
rect 464782 654938 464866 655174
rect 465102 654938 484546 655174
rect 484782 654938 484866 655174
rect 485102 654938 504546 655174
rect 504782 654938 504866 655174
rect 505102 654938 524546 655174
rect 524782 654938 524866 655174
rect 525102 654938 544546 655174
rect 544782 654938 544866 655174
rect 545102 654938 564546 655174
rect 564782 654938 564866 655174
rect 565102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 4546 654854
rect 4782 654618 4866 654854
rect 5102 654618 24546 654854
rect 24782 654618 24866 654854
rect 25102 654618 44546 654854
rect 44782 654618 44866 654854
rect 45102 654618 64546 654854
rect 64782 654618 64866 654854
rect 65102 654618 84546 654854
rect 84782 654618 84866 654854
rect 85102 654618 104546 654854
rect 104782 654618 104866 654854
rect 105102 654618 124546 654854
rect 124782 654618 124866 654854
rect 125102 654618 144546 654854
rect 144782 654618 144866 654854
rect 145102 654618 164546 654854
rect 164782 654618 164866 654854
rect 165102 654618 184546 654854
rect 184782 654618 184866 654854
rect 185102 654618 204546 654854
rect 204782 654618 204866 654854
rect 205102 654618 224546 654854
rect 224782 654618 224866 654854
rect 225102 654618 244546 654854
rect 244782 654618 244866 654854
rect 245102 654618 264546 654854
rect 264782 654618 264866 654854
rect 265102 654618 284546 654854
rect 284782 654618 284866 654854
rect 285102 654618 304546 654854
rect 304782 654618 304866 654854
rect 305102 654618 324546 654854
rect 324782 654618 324866 654854
rect 325102 654618 344546 654854
rect 344782 654618 344866 654854
rect 345102 654618 364546 654854
rect 364782 654618 364866 654854
rect 365102 654618 384546 654854
rect 384782 654618 384866 654854
rect 385102 654618 404546 654854
rect 404782 654618 404866 654854
rect 405102 654618 424546 654854
rect 424782 654618 424866 654854
rect 425102 654618 444546 654854
rect 444782 654618 444866 654854
rect 445102 654618 464546 654854
rect 464782 654618 464866 654854
rect 465102 654618 484546 654854
rect 484782 654618 484866 654854
rect 485102 654618 504546 654854
rect 504782 654618 504866 654854
rect 505102 654618 524546 654854
rect 524782 654618 524866 654854
rect 525102 654618 544546 654854
rect 544782 654618 544866 654854
rect 545102 654618 564546 654854
rect 564782 654618 564866 654854
rect 565102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 826 651454
rect 1062 651218 1146 651454
rect 1382 651218 20826 651454
rect 21062 651218 21146 651454
rect 21382 651218 40826 651454
rect 41062 651218 41146 651454
rect 41382 651218 60826 651454
rect 61062 651218 61146 651454
rect 61382 651218 80826 651454
rect 81062 651218 81146 651454
rect 81382 651218 100826 651454
rect 101062 651218 101146 651454
rect 101382 651218 120826 651454
rect 121062 651218 121146 651454
rect 121382 651218 140826 651454
rect 141062 651218 141146 651454
rect 141382 651218 160826 651454
rect 161062 651218 161146 651454
rect 161382 651218 180826 651454
rect 181062 651218 181146 651454
rect 181382 651218 200826 651454
rect 201062 651218 201146 651454
rect 201382 651218 220826 651454
rect 221062 651218 221146 651454
rect 221382 651218 240826 651454
rect 241062 651218 241146 651454
rect 241382 651218 260826 651454
rect 261062 651218 261146 651454
rect 261382 651218 280826 651454
rect 281062 651218 281146 651454
rect 281382 651218 300826 651454
rect 301062 651218 301146 651454
rect 301382 651218 320826 651454
rect 321062 651218 321146 651454
rect 321382 651218 340826 651454
rect 341062 651218 341146 651454
rect 341382 651218 360826 651454
rect 361062 651218 361146 651454
rect 361382 651218 380826 651454
rect 381062 651218 381146 651454
rect 381382 651218 400826 651454
rect 401062 651218 401146 651454
rect 401382 651218 420826 651454
rect 421062 651218 421146 651454
rect 421382 651218 440826 651454
rect 441062 651218 441146 651454
rect 441382 651218 460826 651454
rect 461062 651218 461146 651454
rect 461382 651218 480826 651454
rect 481062 651218 481146 651454
rect 481382 651218 500826 651454
rect 501062 651218 501146 651454
rect 501382 651218 520826 651454
rect 521062 651218 521146 651454
rect 521382 651218 540826 651454
rect 541062 651218 541146 651454
rect 541382 651218 560826 651454
rect 561062 651218 561146 651454
rect 561382 651218 580826 651454
rect 581062 651218 581146 651454
rect 581382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 826 651134
rect 1062 650898 1146 651134
rect 1382 650898 20826 651134
rect 21062 650898 21146 651134
rect 21382 650898 40826 651134
rect 41062 650898 41146 651134
rect 41382 650898 60826 651134
rect 61062 650898 61146 651134
rect 61382 650898 80826 651134
rect 81062 650898 81146 651134
rect 81382 650898 100826 651134
rect 101062 650898 101146 651134
rect 101382 650898 120826 651134
rect 121062 650898 121146 651134
rect 121382 650898 140826 651134
rect 141062 650898 141146 651134
rect 141382 650898 160826 651134
rect 161062 650898 161146 651134
rect 161382 650898 180826 651134
rect 181062 650898 181146 651134
rect 181382 650898 200826 651134
rect 201062 650898 201146 651134
rect 201382 650898 220826 651134
rect 221062 650898 221146 651134
rect 221382 650898 240826 651134
rect 241062 650898 241146 651134
rect 241382 650898 260826 651134
rect 261062 650898 261146 651134
rect 261382 650898 280826 651134
rect 281062 650898 281146 651134
rect 281382 650898 300826 651134
rect 301062 650898 301146 651134
rect 301382 650898 320826 651134
rect 321062 650898 321146 651134
rect 321382 650898 340826 651134
rect 341062 650898 341146 651134
rect 341382 650898 360826 651134
rect 361062 650898 361146 651134
rect 361382 650898 380826 651134
rect 381062 650898 381146 651134
rect 381382 650898 400826 651134
rect 401062 650898 401146 651134
rect 401382 650898 420826 651134
rect 421062 650898 421146 651134
rect 421382 650898 440826 651134
rect 441062 650898 441146 651134
rect 441382 650898 460826 651134
rect 461062 650898 461146 651134
rect 461382 650898 480826 651134
rect 481062 650898 481146 651134
rect 481382 650898 500826 651134
rect 501062 650898 501146 651134
rect 501382 650898 520826 651134
rect 521062 650898 521146 651134
rect 521382 650898 540826 651134
rect 541062 650898 541146 651134
rect 541382 650898 560826 651134
rect 561062 650898 561146 651134
rect 561382 650898 580826 651134
rect 581062 650898 581146 651134
rect 581382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 21986 644614
rect 22222 644378 22306 644614
rect 22542 644378 41986 644614
rect 42222 644378 42306 644614
rect 42542 644378 61986 644614
rect 62222 644378 62306 644614
rect 62542 644378 81986 644614
rect 82222 644378 82306 644614
rect 82542 644378 101986 644614
rect 102222 644378 102306 644614
rect 102542 644378 121986 644614
rect 122222 644378 122306 644614
rect 122542 644378 141986 644614
rect 142222 644378 142306 644614
rect 142542 644378 161986 644614
rect 162222 644378 162306 644614
rect 162542 644378 181986 644614
rect 182222 644378 182306 644614
rect 182542 644378 201986 644614
rect 202222 644378 202306 644614
rect 202542 644378 221986 644614
rect 222222 644378 222306 644614
rect 222542 644378 241986 644614
rect 242222 644378 242306 644614
rect 242542 644378 261986 644614
rect 262222 644378 262306 644614
rect 262542 644378 281986 644614
rect 282222 644378 282306 644614
rect 282542 644378 301986 644614
rect 302222 644378 302306 644614
rect 302542 644378 321986 644614
rect 322222 644378 322306 644614
rect 322542 644378 341986 644614
rect 342222 644378 342306 644614
rect 342542 644378 361986 644614
rect 362222 644378 362306 644614
rect 362542 644378 381986 644614
rect 382222 644378 382306 644614
rect 382542 644378 401986 644614
rect 402222 644378 402306 644614
rect 402542 644378 421986 644614
rect 422222 644378 422306 644614
rect 422542 644378 441986 644614
rect 442222 644378 442306 644614
rect 442542 644378 461986 644614
rect 462222 644378 462306 644614
rect 462542 644378 481986 644614
rect 482222 644378 482306 644614
rect 482542 644378 501986 644614
rect 502222 644378 502306 644614
rect 502542 644378 521986 644614
rect 522222 644378 522306 644614
rect 522542 644378 541986 644614
rect 542222 644378 542306 644614
rect 542542 644378 561986 644614
rect 562222 644378 562306 644614
rect 562542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 21986 644294
rect 22222 644058 22306 644294
rect 22542 644058 41986 644294
rect 42222 644058 42306 644294
rect 42542 644058 61986 644294
rect 62222 644058 62306 644294
rect 62542 644058 81986 644294
rect 82222 644058 82306 644294
rect 82542 644058 101986 644294
rect 102222 644058 102306 644294
rect 102542 644058 121986 644294
rect 122222 644058 122306 644294
rect 122542 644058 141986 644294
rect 142222 644058 142306 644294
rect 142542 644058 161986 644294
rect 162222 644058 162306 644294
rect 162542 644058 181986 644294
rect 182222 644058 182306 644294
rect 182542 644058 201986 644294
rect 202222 644058 202306 644294
rect 202542 644058 221986 644294
rect 222222 644058 222306 644294
rect 222542 644058 241986 644294
rect 242222 644058 242306 644294
rect 242542 644058 261986 644294
rect 262222 644058 262306 644294
rect 262542 644058 281986 644294
rect 282222 644058 282306 644294
rect 282542 644058 301986 644294
rect 302222 644058 302306 644294
rect 302542 644058 321986 644294
rect 322222 644058 322306 644294
rect 322542 644058 341986 644294
rect 342222 644058 342306 644294
rect 342542 644058 361986 644294
rect 362222 644058 362306 644294
rect 362542 644058 381986 644294
rect 382222 644058 382306 644294
rect 382542 644058 401986 644294
rect 402222 644058 402306 644294
rect 402542 644058 421986 644294
rect 422222 644058 422306 644294
rect 422542 644058 441986 644294
rect 442222 644058 442306 644294
rect 442542 644058 461986 644294
rect 462222 644058 462306 644294
rect 462542 644058 481986 644294
rect 482222 644058 482306 644294
rect 482542 644058 501986 644294
rect 502222 644058 502306 644294
rect 502542 644058 521986 644294
rect 522222 644058 522306 644294
rect 522542 644058 541986 644294
rect 542222 644058 542306 644294
rect 542542 644058 561986 644294
rect 562222 644058 562306 644294
rect 562542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 18266 640894
rect 18502 640658 18586 640894
rect 18822 640658 38266 640894
rect 38502 640658 38586 640894
rect 38822 640658 58266 640894
rect 58502 640658 58586 640894
rect 58822 640658 78266 640894
rect 78502 640658 78586 640894
rect 78822 640658 98266 640894
rect 98502 640658 98586 640894
rect 98822 640658 118266 640894
rect 118502 640658 118586 640894
rect 118822 640658 138266 640894
rect 138502 640658 138586 640894
rect 138822 640658 158266 640894
rect 158502 640658 158586 640894
rect 158822 640658 178266 640894
rect 178502 640658 178586 640894
rect 178822 640658 198266 640894
rect 198502 640658 198586 640894
rect 198822 640658 218266 640894
rect 218502 640658 218586 640894
rect 218822 640658 238266 640894
rect 238502 640658 238586 640894
rect 238822 640658 258266 640894
rect 258502 640658 258586 640894
rect 258822 640658 278266 640894
rect 278502 640658 278586 640894
rect 278822 640658 298266 640894
rect 298502 640658 298586 640894
rect 298822 640658 318266 640894
rect 318502 640658 318586 640894
rect 318822 640658 338266 640894
rect 338502 640658 338586 640894
rect 338822 640658 358266 640894
rect 358502 640658 358586 640894
rect 358822 640658 378266 640894
rect 378502 640658 378586 640894
rect 378822 640658 398266 640894
rect 398502 640658 398586 640894
rect 398822 640658 418266 640894
rect 418502 640658 418586 640894
rect 418822 640658 438266 640894
rect 438502 640658 438586 640894
rect 438822 640658 458266 640894
rect 458502 640658 458586 640894
rect 458822 640658 478266 640894
rect 478502 640658 478586 640894
rect 478822 640658 498266 640894
rect 498502 640658 498586 640894
rect 498822 640658 518266 640894
rect 518502 640658 518586 640894
rect 518822 640658 538266 640894
rect 538502 640658 538586 640894
rect 538822 640658 558266 640894
rect 558502 640658 558586 640894
rect 558822 640658 578266 640894
rect 578502 640658 578586 640894
rect 578822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 18266 640574
rect 18502 640338 18586 640574
rect 18822 640338 38266 640574
rect 38502 640338 38586 640574
rect 38822 640338 58266 640574
rect 58502 640338 58586 640574
rect 58822 640338 78266 640574
rect 78502 640338 78586 640574
rect 78822 640338 98266 640574
rect 98502 640338 98586 640574
rect 98822 640338 118266 640574
rect 118502 640338 118586 640574
rect 118822 640338 138266 640574
rect 138502 640338 138586 640574
rect 138822 640338 158266 640574
rect 158502 640338 158586 640574
rect 158822 640338 178266 640574
rect 178502 640338 178586 640574
rect 178822 640338 198266 640574
rect 198502 640338 198586 640574
rect 198822 640338 218266 640574
rect 218502 640338 218586 640574
rect 218822 640338 238266 640574
rect 238502 640338 238586 640574
rect 238822 640338 258266 640574
rect 258502 640338 258586 640574
rect 258822 640338 278266 640574
rect 278502 640338 278586 640574
rect 278822 640338 298266 640574
rect 298502 640338 298586 640574
rect 298822 640338 318266 640574
rect 318502 640338 318586 640574
rect 318822 640338 338266 640574
rect 338502 640338 338586 640574
rect 338822 640338 358266 640574
rect 358502 640338 358586 640574
rect 358822 640338 378266 640574
rect 378502 640338 378586 640574
rect 378822 640338 398266 640574
rect 398502 640338 398586 640574
rect 398822 640338 418266 640574
rect 418502 640338 418586 640574
rect 418822 640338 438266 640574
rect 438502 640338 438586 640574
rect 438822 640338 458266 640574
rect 458502 640338 458586 640574
rect 458822 640338 478266 640574
rect 478502 640338 478586 640574
rect 478822 640338 498266 640574
rect 498502 640338 498586 640574
rect 498822 640338 518266 640574
rect 518502 640338 518586 640574
rect 518822 640338 538266 640574
rect 538502 640338 538586 640574
rect 538822 640338 558266 640574
rect 558502 640338 558586 640574
rect 558822 640338 578266 640574
rect 578502 640338 578586 640574
rect 578822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 14546 637174
rect 14782 636938 14866 637174
rect 15102 636938 34546 637174
rect 34782 636938 34866 637174
rect 35102 636938 54546 637174
rect 54782 636938 54866 637174
rect 55102 636938 74546 637174
rect 74782 636938 74866 637174
rect 75102 636938 94546 637174
rect 94782 636938 94866 637174
rect 95102 636938 114546 637174
rect 114782 636938 114866 637174
rect 115102 636938 134546 637174
rect 134782 636938 134866 637174
rect 135102 636938 154546 637174
rect 154782 636938 154866 637174
rect 155102 636938 174546 637174
rect 174782 636938 174866 637174
rect 175102 636938 194546 637174
rect 194782 636938 194866 637174
rect 195102 636938 214546 637174
rect 214782 636938 214866 637174
rect 215102 636938 234546 637174
rect 234782 636938 234866 637174
rect 235102 636938 254546 637174
rect 254782 636938 254866 637174
rect 255102 636938 274546 637174
rect 274782 636938 274866 637174
rect 275102 636938 294546 637174
rect 294782 636938 294866 637174
rect 295102 636938 314546 637174
rect 314782 636938 314866 637174
rect 315102 636938 334546 637174
rect 334782 636938 334866 637174
rect 335102 636938 354546 637174
rect 354782 636938 354866 637174
rect 355102 636938 374546 637174
rect 374782 636938 374866 637174
rect 375102 636938 394546 637174
rect 394782 636938 394866 637174
rect 395102 636938 414546 637174
rect 414782 636938 414866 637174
rect 415102 636938 434546 637174
rect 434782 636938 434866 637174
rect 435102 636938 454546 637174
rect 454782 636938 454866 637174
rect 455102 636938 474546 637174
rect 474782 636938 474866 637174
rect 475102 636938 494546 637174
rect 494782 636938 494866 637174
rect 495102 636938 514546 637174
rect 514782 636938 514866 637174
rect 515102 636938 534546 637174
rect 534782 636938 534866 637174
rect 535102 636938 554546 637174
rect 554782 636938 554866 637174
rect 555102 636938 574546 637174
rect 574782 636938 574866 637174
rect 575102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 14546 636854
rect 14782 636618 14866 636854
rect 15102 636618 34546 636854
rect 34782 636618 34866 636854
rect 35102 636618 54546 636854
rect 54782 636618 54866 636854
rect 55102 636618 74546 636854
rect 74782 636618 74866 636854
rect 75102 636618 94546 636854
rect 94782 636618 94866 636854
rect 95102 636618 114546 636854
rect 114782 636618 114866 636854
rect 115102 636618 134546 636854
rect 134782 636618 134866 636854
rect 135102 636618 154546 636854
rect 154782 636618 154866 636854
rect 155102 636618 174546 636854
rect 174782 636618 174866 636854
rect 175102 636618 194546 636854
rect 194782 636618 194866 636854
rect 195102 636618 214546 636854
rect 214782 636618 214866 636854
rect 215102 636618 234546 636854
rect 234782 636618 234866 636854
rect 235102 636618 254546 636854
rect 254782 636618 254866 636854
rect 255102 636618 274546 636854
rect 274782 636618 274866 636854
rect 275102 636618 294546 636854
rect 294782 636618 294866 636854
rect 295102 636618 314546 636854
rect 314782 636618 314866 636854
rect 315102 636618 334546 636854
rect 334782 636618 334866 636854
rect 335102 636618 354546 636854
rect 354782 636618 354866 636854
rect 355102 636618 374546 636854
rect 374782 636618 374866 636854
rect 375102 636618 394546 636854
rect 394782 636618 394866 636854
rect 395102 636618 414546 636854
rect 414782 636618 414866 636854
rect 415102 636618 434546 636854
rect 434782 636618 434866 636854
rect 435102 636618 454546 636854
rect 454782 636618 454866 636854
rect 455102 636618 474546 636854
rect 474782 636618 474866 636854
rect 475102 636618 494546 636854
rect 494782 636618 494866 636854
rect 495102 636618 514546 636854
rect 514782 636618 514866 636854
rect 515102 636618 534546 636854
rect 534782 636618 534866 636854
rect 535102 636618 554546 636854
rect 554782 636618 554866 636854
rect 555102 636618 574546 636854
rect 574782 636618 574866 636854
rect 575102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 10826 633454
rect 11062 633218 11146 633454
rect 11382 633218 30826 633454
rect 31062 633218 31146 633454
rect 31382 633218 50826 633454
rect 51062 633218 51146 633454
rect 51382 633218 70826 633454
rect 71062 633218 71146 633454
rect 71382 633218 90826 633454
rect 91062 633218 91146 633454
rect 91382 633218 110826 633454
rect 111062 633218 111146 633454
rect 111382 633218 130826 633454
rect 131062 633218 131146 633454
rect 131382 633218 150826 633454
rect 151062 633218 151146 633454
rect 151382 633218 170826 633454
rect 171062 633218 171146 633454
rect 171382 633218 190826 633454
rect 191062 633218 191146 633454
rect 191382 633218 210826 633454
rect 211062 633218 211146 633454
rect 211382 633218 230826 633454
rect 231062 633218 231146 633454
rect 231382 633218 250826 633454
rect 251062 633218 251146 633454
rect 251382 633218 270826 633454
rect 271062 633218 271146 633454
rect 271382 633218 290826 633454
rect 291062 633218 291146 633454
rect 291382 633218 310826 633454
rect 311062 633218 311146 633454
rect 311382 633218 330826 633454
rect 331062 633218 331146 633454
rect 331382 633218 350826 633454
rect 351062 633218 351146 633454
rect 351382 633218 370826 633454
rect 371062 633218 371146 633454
rect 371382 633218 390826 633454
rect 391062 633218 391146 633454
rect 391382 633218 410826 633454
rect 411062 633218 411146 633454
rect 411382 633218 430826 633454
rect 431062 633218 431146 633454
rect 431382 633218 450826 633454
rect 451062 633218 451146 633454
rect 451382 633218 470826 633454
rect 471062 633218 471146 633454
rect 471382 633218 490826 633454
rect 491062 633218 491146 633454
rect 491382 633218 510826 633454
rect 511062 633218 511146 633454
rect 511382 633218 530826 633454
rect 531062 633218 531146 633454
rect 531382 633218 550826 633454
rect 551062 633218 551146 633454
rect 551382 633218 570826 633454
rect 571062 633218 571146 633454
rect 571382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 10826 633134
rect 11062 632898 11146 633134
rect 11382 632898 30826 633134
rect 31062 632898 31146 633134
rect 31382 632898 50826 633134
rect 51062 632898 51146 633134
rect 51382 632898 70826 633134
rect 71062 632898 71146 633134
rect 71382 632898 90826 633134
rect 91062 632898 91146 633134
rect 91382 632898 110826 633134
rect 111062 632898 111146 633134
rect 111382 632898 130826 633134
rect 131062 632898 131146 633134
rect 131382 632898 150826 633134
rect 151062 632898 151146 633134
rect 151382 632898 170826 633134
rect 171062 632898 171146 633134
rect 171382 632898 190826 633134
rect 191062 632898 191146 633134
rect 191382 632898 210826 633134
rect 211062 632898 211146 633134
rect 211382 632898 230826 633134
rect 231062 632898 231146 633134
rect 231382 632898 250826 633134
rect 251062 632898 251146 633134
rect 251382 632898 270826 633134
rect 271062 632898 271146 633134
rect 271382 632898 290826 633134
rect 291062 632898 291146 633134
rect 291382 632898 310826 633134
rect 311062 632898 311146 633134
rect 311382 632898 330826 633134
rect 331062 632898 331146 633134
rect 331382 632898 350826 633134
rect 351062 632898 351146 633134
rect 351382 632898 370826 633134
rect 371062 632898 371146 633134
rect 371382 632898 390826 633134
rect 391062 632898 391146 633134
rect 391382 632898 410826 633134
rect 411062 632898 411146 633134
rect 411382 632898 430826 633134
rect 431062 632898 431146 633134
rect 431382 632898 450826 633134
rect 451062 632898 451146 633134
rect 451382 632898 470826 633134
rect 471062 632898 471146 633134
rect 471382 632898 490826 633134
rect 491062 632898 491146 633134
rect 491382 632898 510826 633134
rect 511062 632898 511146 633134
rect 511382 632898 530826 633134
rect 531062 632898 531146 633134
rect 531382 632898 550826 633134
rect 551062 632898 551146 633134
rect 551382 632898 570826 633134
rect 571062 632898 571146 633134
rect 571382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 11986 626614
rect 12222 626378 12306 626614
rect 12542 626378 31986 626614
rect 32222 626378 32306 626614
rect 32542 626378 51986 626614
rect 52222 626378 52306 626614
rect 52542 626378 71986 626614
rect 72222 626378 72306 626614
rect 72542 626378 91986 626614
rect 92222 626378 92306 626614
rect 92542 626378 111986 626614
rect 112222 626378 112306 626614
rect 112542 626378 131986 626614
rect 132222 626378 132306 626614
rect 132542 626378 151986 626614
rect 152222 626378 152306 626614
rect 152542 626378 171986 626614
rect 172222 626378 172306 626614
rect 172542 626378 191986 626614
rect 192222 626378 192306 626614
rect 192542 626378 211986 626614
rect 212222 626378 212306 626614
rect 212542 626378 231986 626614
rect 232222 626378 232306 626614
rect 232542 626378 251986 626614
rect 252222 626378 252306 626614
rect 252542 626378 271986 626614
rect 272222 626378 272306 626614
rect 272542 626378 291986 626614
rect 292222 626378 292306 626614
rect 292542 626378 311986 626614
rect 312222 626378 312306 626614
rect 312542 626378 331986 626614
rect 332222 626378 332306 626614
rect 332542 626378 351986 626614
rect 352222 626378 352306 626614
rect 352542 626378 371986 626614
rect 372222 626378 372306 626614
rect 372542 626378 391986 626614
rect 392222 626378 392306 626614
rect 392542 626378 411986 626614
rect 412222 626378 412306 626614
rect 412542 626378 431986 626614
rect 432222 626378 432306 626614
rect 432542 626378 451986 626614
rect 452222 626378 452306 626614
rect 452542 626378 471986 626614
rect 472222 626378 472306 626614
rect 472542 626378 491986 626614
rect 492222 626378 492306 626614
rect 492542 626378 511986 626614
rect 512222 626378 512306 626614
rect 512542 626378 531986 626614
rect 532222 626378 532306 626614
rect 532542 626378 551986 626614
rect 552222 626378 552306 626614
rect 552542 626378 571986 626614
rect 572222 626378 572306 626614
rect 572542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 11986 626294
rect 12222 626058 12306 626294
rect 12542 626058 31986 626294
rect 32222 626058 32306 626294
rect 32542 626058 51986 626294
rect 52222 626058 52306 626294
rect 52542 626058 71986 626294
rect 72222 626058 72306 626294
rect 72542 626058 91986 626294
rect 92222 626058 92306 626294
rect 92542 626058 111986 626294
rect 112222 626058 112306 626294
rect 112542 626058 131986 626294
rect 132222 626058 132306 626294
rect 132542 626058 151986 626294
rect 152222 626058 152306 626294
rect 152542 626058 171986 626294
rect 172222 626058 172306 626294
rect 172542 626058 191986 626294
rect 192222 626058 192306 626294
rect 192542 626058 211986 626294
rect 212222 626058 212306 626294
rect 212542 626058 231986 626294
rect 232222 626058 232306 626294
rect 232542 626058 251986 626294
rect 252222 626058 252306 626294
rect 252542 626058 271986 626294
rect 272222 626058 272306 626294
rect 272542 626058 291986 626294
rect 292222 626058 292306 626294
rect 292542 626058 311986 626294
rect 312222 626058 312306 626294
rect 312542 626058 331986 626294
rect 332222 626058 332306 626294
rect 332542 626058 351986 626294
rect 352222 626058 352306 626294
rect 352542 626058 371986 626294
rect 372222 626058 372306 626294
rect 372542 626058 391986 626294
rect 392222 626058 392306 626294
rect 392542 626058 411986 626294
rect 412222 626058 412306 626294
rect 412542 626058 431986 626294
rect 432222 626058 432306 626294
rect 432542 626058 451986 626294
rect 452222 626058 452306 626294
rect 452542 626058 471986 626294
rect 472222 626058 472306 626294
rect 472542 626058 491986 626294
rect 492222 626058 492306 626294
rect 492542 626058 511986 626294
rect 512222 626058 512306 626294
rect 512542 626058 531986 626294
rect 532222 626058 532306 626294
rect 532542 626058 551986 626294
rect 552222 626058 552306 626294
rect 552542 626058 571986 626294
rect 572222 626058 572306 626294
rect 572542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 8266 622894
rect 8502 622658 8586 622894
rect 8822 622658 28266 622894
rect 28502 622658 28586 622894
rect 28822 622658 48266 622894
rect 48502 622658 48586 622894
rect 48822 622658 68266 622894
rect 68502 622658 68586 622894
rect 68822 622658 88266 622894
rect 88502 622658 88586 622894
rect 88822 622658 108266 622894
rect 108502 622658 108586 622894
rect 108822 622658 128266 622894
rect 128502 622658 128586 622894
rect 128822 622658 148266 622894
rect 148502 622658 148586 622894
rect 148822 622658 168266 622894
rect 168502 622658 168586 622894
rect 168822 622658 188266 622894
rect 188502 622658 188586 622894
rect 188822 622658 208266 622894
rect 208502 622658 208586 622894
rect 208822 622658 228266 622894
rect 228502 622658 228586 622894
rect 228822 622658 248266 622894
rect 248502 622658 248586 622894
rect 248822 622658 268266 622894
rect 268502 622658 268586 622894
rect 268822 622658 288266 622894
rect 288502 622658 288586 622894
rect 288822 622658 308266 622894
rect 308502 622658 308586 622894
rect 308822 622658 328266 622894
rect 328502 622658 328586 622894
rect 328822 622658 348266 622894
rect 348502 622658 348586 622894
rect 348822 622658 368266 622894
rect 368502 622658 368586 622894
rect 368822 622658 388266 622894
rect 388502 622658 388586 622894
rect 388822 622658 408266 622894
rect 408502 622658 408586 622894
rect 408822 622658 428266 622894
rect 428502 622658 428586 622894
rect 428822 622658 448266 622894
rect 448502 622658 448586 622894
rect 448822 622658 468266 622894
rect 468502 622658 468586 622894
rect 468822 622658 488266 622894
rect 488502 622658 488586 622894
rect 488822 622658 508266 622894
rect 508502 622658 508586 622894
rect 508822 622658 528266 622894
rect 528502 622658 528586 622894
rect 528822 622658 548266 622894
rect 548502 622658 548586 622894
rect 548822 622658 568266 622894
rect 568502 622658 568586 622894
rect 568822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 8266 622574
rect 8502 622338 8586 622574
rect 8822 622338 28266 622574
rect 28502 622338 28586 622574
rect 28822 622338 48266 622574
rect 48502 622338 48586 622574
rect 48822 622338 68266 622574
rect 68502 622338 68586 622574
rect 68822 622338 88266 622574
rect 88502 622338 88586 622574
rect 88822 622338 108266 622574
rect 108502 622338 108586 622574
rect 108822 622338 128266 622574
rect 128502 622338 128586 622574
rect 128822 622338 148266 622574
rect 148502 622338 148586 622574
rect 148822 622338 168266 622574
rect 168502 622338 168586 622574
rect 168822 622338 188266 622574
rect 188502 622338 188586 622574
rect 188822 622338 208266 622574
rect 208502 622338 208586 622574
rect 208822 622338 228266 622574
rect 228502 622338 228586 622574
rect 228822 622338 248266 622574
rect 248502 622338 248586 622574
rect 248822 622338 268266 622574
rect 268502 622338 268586 622574
rect 268822 622338 288266 622574
rect 288502 622338 288586 622574
rect 288822 622338 308266 622574
rect 308502 622338 308586 622574
rect 308822 622338 328266 622574
rect 328502 622338 328586 622574
rect 328822 622338 348266 622574
rect 348502 622338 348586 622574
rect 348822 622338 368266 622574
rect 368502 622338 368586 622574
rect 368822 622338 388266 622574
rect 388502 622338 388586 622574
rect 388822 622338 408266 622574
rect 408502 622338 408586 622574
rect 408822 622338 428266 622574
rect 428502 622338 428586 622574
rect 428822 622338 448266 622574
rect 448502 622338 448586 622574
rect 448822 622338 468266 622574
rect 468502 622338 468586 622574
rect 468822 622338 488266 622574
rect 488502 622338 488586 622574
rect 488822 622338 508266 622574
rect 508502 622338 508586 622574
rect 508822 622338 528266 622574
rect 528502 622338 528586 622574
rect 528822 622338 548266 622574
rect 548502 622338 548586 622574
rect 548822 622338 568266 622574
rect 568502 622338 568586 622574
rect 568822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 4546 619174
rect 4782 618938 4866 619174
rect 5102 618938 24546 619174
rect 24782 618938 24866 619174
rect 25102 618938 44546 619174
rect 44782 618938 44866 619174
rect 45102 618938 64546 619174
rect 64782 618938 64866 619174
rect 65102 618938 84546 619174
rect 84782 618938 84866 619174
rect 85102 618938 104546 619174
rect 104782 618938 104866 619174
rect 105102 618938 124546 619174
rect 124782 618938 124866 619174
rect 125102 618938 144546 619174
rect 144782 618938 144866 619174
rect 145102 618938 164546 619174
rect 164782 618938 164866 619174
rect 165102 618938 184546 619174
rect 184782 618938 184866 619174
rect 185102 618938 204546 619174
rect 204782 618938 204866 619174
rect 205102 618938 224546 619174
rect 224782 618938 224866 619174
rect 225102 618938 244546 619174
rect 244782 618938 244866 619174
rect 245102 618938 264546 619174
rect 264782 618938 264866 619174
rect 265102 618938 284546 619174
rect 284782 618938 284866 619174
rect 285102 618938 304546 619174
rect 304782 618938 304866 619174
rect 305102 618938 324546 619174
rect 324782 618938 324866 619174
rect 325102 618938 344546 619174
rect 344782 618938 344866 619174
rect 345102 618938 364546 619174
rect 364782 618938 364866 619174
rect 365102 618938 384546 619174
rect 384782 618938 384866 619174
rect 385102 618938 404546 619174
rect 404782 618938 404866 619174
rect 405102 618938 424546 619174
rect 424782 618938 424866 619174
rect 425102 618938 444546 619174
rect 444782 618938 444866 619174
rect 445102 618938 464546 619174
rect 464782 618938 464866 619174
rect 465102 618938 484546 619174
rect 484782 618938 484866 619174
rect 485102 618938 504546 619174
rect 504782 618938 504866 619174
rect 505102 618938 524546 619174
rect 524782 618938 524866 619174
rect 525102 618938 544546 619174
rect 544782 618938 544866 619174
rect 545102 618938 564546 619174
rect 564782 618938 564866 619174
rect 565102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 4546 618854
rect 4782 618618 4866 618854
rect 5102 618618 24546 618854
rect 24782 618618 24866 618854
rect 25102 618618 44546 618854
rect 44782 618618 44866 618854
rect 45102 618618 64546 618854
rect 64782 618618 64866 618854
rect 65102 618618 84546 618854
rect 84782 618618 84866 618854
rect 85102 618618 104546 618854
rect 104782 618618 104866 618854
rect 105102 618618 124546 618854
rect 124782 618618 124866 618854
rect 125102 618618 144546 618854
rect 144782 618618 144866 618854
rect 145102 618618 164546 618854
rect 164782 618618 164866 618854
rect 165102 618618 184546 618854
rect 184782 618618 184866 618854
rect 185102 618618 204546 618854
rect 204782 618618 204866 618854
rect 205102 618618 224546 618854
rect 224782 618618 224866 618854
rect 225102 618618 244546 618854
rect 244782 618618 244866 618854
rect 245102 618618 264546 618854
rect 264782 618618 264866 618854
rect 265102 618618 284546 618854
rect 284782 618618 284866 618854
rect 285102 618618 304546 618854
rect 304782 618618 304866 618854
rect 305102 618618 324546 618854
rect 324782 618618 324866 618854
rect 325102 618618 344546 618854
rect 344782 618618 344866 618854
rect 345102 618618 364546 618854
rect 364782 618618 364866 618854
rect 365102 618618 384546 618854
rect 384782 618618 384866 618854
rect 385102 618618 404546 618854
rect 404782 618618 404866 618854
rect 405102 618618 424546 618854
rect 424782 618618 424866 618854
rect 425102 618618 444546 618854
rect 444782 618618 444866 618854
rect 445102 618618 464546 618854
rect 464782 618618 464866 618854
rect 465102 618618 484546 618854
rect 484782 618618 484866 618854
rect 485102 618618 504546 618854
rect 504782 618618 504866 618854
rect 505102 618618 524546 618854
rect 524782 618618 524866 618854
rect 525102 618618 544546 618854
rect 544782 618618 544866 618854
rect 545102 618618 564546 618854
rect 564782 618618 564866 618854
rect 565102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 826 615454
rect 1062 615218 1146 615454
rect 1382 615218 20826 615454
rect 21062 615218 21146 615454
rect 21382 615218 40826 615454
rect 41062 615218 41146 615454
rect 41382 615218 60826 615454
rect 61062 615218 61146 615454
rect 61382 615218 80826 615454
rect 81062 615218 81146 615454
rect 81382 615218 100826 615454
rect 101062 615218 101146 615454
rect 101382 615218 120826 615454
rect 121062 615218 121146 615454
rect 121382 615218 140826 615454
rect 141062 615218 141146 615454
rect 141382 615218 160826 615454
rect 161062 615218 161146 615454
rect 161382 615218 180826 615454
rect 181062 615218 181146 615454
rect 181382 615218 200826 615454
rect 201062 615218 201146 615454
rect 201382 615218 220826 615454
rect 221062 615218 221146 615454
rect 221382 615218 240826 615454
rect 241062 615218 241146 615454
rect 241382 615218 260826 615454
rect 261062 615218 261146 615454
rect 261382 615218 280826 615454
rect 281062 615218 281146 615454
rect 281382 615218 300826 615454
rect 301062 615218 301146 615454
rect 301382 615218 320826 615454
rect 321062 615218 321146 615454
rect 321382 615218 340826 615454
rect 341062 615218 341146 615454
rect 341382 615218 360826 615454
rect 361062 615218 361146 615454
rect 361382 615218 380826 615454
rect 381062 615218 381146 615454
rect 381382 615218 400826 615454
rect 401062 615218 401146 615454
rect 401382 615218 420826 615454
rect 421062 615218 421146 615454
rect 421382 615218 440826 615454
rect 441062 615218 441146 615454
rect 441382 615218 460826 615454
rect 461062 615218 461146 615454
rect 461382 615218 480826 615454
rect 481062 615218 481146 615454
rect 481382 615218 500826 615454
rect 501062 615218 501146 615454
rect 501382 615218 520826 615454
rect 521062 615218 521146 615454
rect 521382 615218 540826 615454
rect 541062 615218 541146 615454
rect 541382 615218 560826 615454
rect 561062 615218 561146 615454
rect 561382 615218 580826 615454
rect 581062 615218 581146 615454
rect 581382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 826 615134
rect 1062 614898 1146 615134
rect 1382 614898 20826 615134
rect 21062 614898 21146 615134
rect 21382 614898 40826 615134
rect 41062 614898 41146 615134
rect 41382 614898 60826 615134
rect 61062 614898 61146 615134
rect 61382 614898 80826 615134
rect 81062 614898 81146 615134
rect 81382 614898 100826 615134
rect 101062 614898 101146 615134
rect 101382 614898 120826 615134
rect 121062 614898 121146 615134
rect 121382 614898 140826 615134
rect 141062 614898 141146 615134
rect 141382 614898 160826 615134
rect 161062 614898 161146 615134
rect 161382 614898 180826 615134
rect 181062 614898 181146 615134
rect 181382 614898 200826 615134
rect 201062 614898 201146 615134
rect 201382 614898 220826 615134
rect 221062 614898 221146 615134
rect 221382 614898 240826 615134
rect 241062 614898 241146 615134
rect 241382 614898 260826 615134
rect 261062 614898 261146 615134
rect 261382 614898 280826 615134
rect 281062 614898 281146 615134
rect 281382 614898 300826 615134
rect 301062 614898 301146 615134
rect 301382 614898 320826 615134
rect 321062 614898 321146 615134
rect 321382 614898 340826 615134
rect 341062 614898 341146 615134
rect 341382 614898 360826 615134
rect 361062 614898 361146 615134
rect 361382 614898 380826 615134
rect 381062 614898 381146 615134
rect 381382 614898 400826 615134
rect 401062 614898 401146 615134
rect 401382 614898 420826 615134
rect 421062 614898 421146 615134
rect 421382 614898 440826 615134
rect 441062 614898 441146 615134
rect 441382 614898 460826 615134
rect 461062 614898 461146 615134
rect 461382 614898 480826 615134
rect 481062 614898 481146 615134
rect 481382 614898 500826 615134
rect 501062 614898 501146 615134
rect 501382 614898 520826 615134
rect 521062 614898 521146 615134
rect 521382 614898 540826 615134
rect 541062 614898 541146 615134
rect 541382 614898 560826 615134
rect 561062 614898 561146 615134
rect 561382 614898 580826 615134
rect 581062 614898 581146 615134
rect 581382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 21986 608614
rect 22222 608378 22306 608614
rect 22542 608378 41986 608614
rect 42222 608378 42306 608614
rect 42542 608378 61986 608614
rect 62222 608378 62306 608614
rect 62542 608378 81986 608614
rect 82222 608378 82306 608614
rect 82542 608378 101986 608614
rect 102222 608378 102306 608614
rect 102542 608378 121986 608614
rect 122222 608378 122306 608614
rect 122542 608378 141986 608614
rect 142222 608378 142306 608614
rect 142542 608378 161986 608614
rect 162222 608378 162306 608614
rect 162542 608378 181986 608614
rect 182222 608378 182306 608614
rect 182542 608378 201986 608614
rect 202222 608378 202306 608614
rect 202542 608378 221986 608614
rect 222222 608378 222306 608614
rect 222542 608378 241986 608614
rect 242222 608378 242306 608614
rect 242542 608378 261986 608614
rect 262222 608378 262306 608614
rect 262542 608378 281986 608614
rect 282222 608378 282306 608614
rect 282542 608378 301986 608614
rect 302222 608378 302306 608614
rect 302542 608378 321986 608614
rect 322222 608378 322306 608614
rect 322542 608378 341986 608614
rect 342222 608378 342306 608614
rect 342542 608378 361986 608614
rect 362222 608378 362306 608614
rect 362542 608378 381986 608614
rect 382222 608378 382306 608614
rect 382542 608378 401986 608614
rect 402222 608378 402306 608614
rect 402542 608378 421986 608614
rect 422222 608378 422306 608614
rect 422542 608378 441986 608614
rect 442222 608378 442306 608614
rect 442542 608378 461986 608614
rect 462222 608378 462306 608614
rect 462542 608378 481986 608614
rect 482222 608378 482306 608614
rect 482542 608378 501986 608614
rect 502222 608378 502306 608614
rect 502542 608378 521986 608614
rect 522222 608378 522306 608614
rect 522542 608378 541986 608614
rect 542222 608378 542306 608614
rect 542542 608378 561986 608614
rect 562222 608378 562306 608614
rect 562542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 21986 608294
rect 22222 608058 22306 608294
rect 22542 608058 41986 608294
rect 42222 608058 42306 608294
rect 42542 608058 61986 608294
rect 62222 608058 62306 608294
rect 62542 608058 81986 608294
rect 82222 608058 82306 608294
rect 82542 608058 101986 608294
rect 102222 608058 102306 608294
rect 102542 608058 121986 608294
rect 122222 608058 122306 608294
rect 122542 608058 141986 608294
rect 142222 608058 142306 608294
rect 142542 608058 161986 608294
rect 162222 608058 162306 608294
rect 162542 608058 181986 608294
rect 182222 608058 182306 608294
rect 182542 608058 201986 608294
rect 202222 608058 202306 608294
rect 202542 608058 221986 608294
rect 222222 608058 222306 608294
rect 222542 608058 241986 608294
rect 242222 608058 242306 608294
rect 242542 608058 261986 608294
rect 262222 608058 262306 608294
rect 262542 608058 281986 608294
rect 282222 608058 282306 608294
rect 282542 608058 301986 608294
rect 302222 608058 302306 608294
rect 302542 608058 321986 608294
rect 322222 608058 322306 608294
rect 322542 608058 341986 608294
rect 342222 608058 342306 608294
rect 342542 608058 361986 608294
rect 362222 608058 362306 608294
rect 362542 608058 381986 608294
rect 382222 608058 382306 608294
rect 382542 608058 401986 608294
rect 402222 608058 402306 608294
rect 402542 608058 421986 608294
rect 422222 608058 422306 608294
rect 422542 608058 441986 608294
rect 442222 608058 442306 608294
rect 442542 608058 461986 608294
rect 462222 608058 462306 608294
rect 462542 608058 481986 608294
rect 482222 608058 482306 608294
rect 482542 608058 501986 608294
rect 502222 608058 502306 608294
rect 502542 608058 521986 608294
rect 522222 608058 522306 608294
rect 522542 608058 541986 608294
rect 542222 608058 542306 608294
rect 542542 608058 561986 608294
rect 562222 608058 562306 608294
rect 562542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 18266 604894
rect 18502 604658 18586 604894
rect 18822 604658 38266 604894
rect 38502 604658 38586 604894
rect 38822 604658 58266 604894
rect 58502 604658 58586 604894
rect 58822 604658 78266 604894
rect 78502 604658 78586 604894
rect 78822 604658 98266 604894
rect 98502 604658 98586 604894
rect 98822 604658 118266 604894
rect 118502 604658 118586 604894
rect 118822 604658 138266 604894
rect 138502 604658 138586 604894
rect 138822 604658 158266 604894
rect 158502 604658 158586 604894
rect 158822 604658 178266 604894
rect 178502 604658 178586 604894
rect 178822 604658 198266 604894
rect 198502 604658 198586 604894
rect 198822 604658 218266 604894
rect 218502 604658 218586 604894
rect 218822 604658 238266 604894
rect 238502 604658 238586 604894
rect 238822 604658 258266 604894
rect 258502 604658 258586 604894
rect 258822 604658 278266 604894
rect 278502 604658 278586 604894
rect 278822 604658 298266 604894
rect 298502 604658 298586 604894
rect 298822 604658 318266 604894
rect 318502 604658 318586 604894
rect 318822 604658 338266 604894
rect 338502 604658 338586 604894
rect 338822 604658 358266 604894
rect 358502 604658 358586 604894
rect 358822 604658 378266 604894
rect 378502 604658 378586 604894
rect 378822 604658 398266 604894
rect 398502 604658 398586 604894
rect 398822 604658 418266 604894
rect 418502 604658 418586 604894
rect 418822 604658 438266 604894
rect 438502 604658 438586 604894
rect 438822 604658 458266 604894
rect 458502 604658 458586 604894
rect 458822 604658 478266 604894
rect 478502 604658 478586 604894
rect 478822 604658 498266 604894
rect 498502 604658 498586 604894
rect 498822 604658 518266 604894
rect 518502 604658 518586 604894
rect 518822 604658 538266 604894
rect 538502 604658 538586 604894
rect 538822 604658 558266 604894
rect 558502 604658 558586 604894
rect 558822 604658 578266 604894
rect 578502 604658 578586 604894
rect 578822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 18266 604574
rect 18502 604338 18586 604574
rect 18822 604338 38266 604574
rect 38502 604338 38586 604574
rect 38822 604338 58266 604574
rect 58502 604338 58586 604574
rect 58822 604338 78266 604574
rect 78502 604338 78586 604574
rect 78822 604338 98266 604574
rect 98502 604338 98586 604574
rect 98822 604338 118266 604574
rect 118502 604338 118586 604574
rect 118822 604338 138266 604574
rect 138502 604338 138586 604574
rect 138822 604338 158266 604574
rect 158502 604338 158586 604574
rect 158822 604338 178266 604574
rect 178502 604338 178586 604574
rect 178822 604338 198266 604574
rect 198502 604338 198586 604574
rect 198822 604338 218266 604574
rect 218502 604338 218586 604574
rect 218822 604338 238266 604574
rect 238502 604338 238586 604574
rect 238822 604338 258266 604574
rect 258502 604338 258586 604574
rect 258822 604338 278266 604574
rect 278502 604338 278586 604574
rect 278822 604338 298266 604574
rect 298502 604338 298586 604574
rect 298822 604338 318266 604574
rect 318502 604338 318586 604574
rect 318822 604338 338266 604574
rect 338502 604338 338586 604574
rect 338822 604338 358266 604574
rect 358502 604338 358586 604574
rect 358822 604338 378266 604574
rect 378502 604338 378586 604574
rect 378822 604338 398266 604574
rect 398502 604338 398586 604574
rect 398822 604338 418266 604574
rect 418502 604338 418586 604574
rect 418822 604338 438266 604574
rect 438502 604338 438586 604574
rect 438822 604338 458266 604574
rect 458502 604338 458586 604574
rect 458822 604338 478266 604574
rect 478502 604338 478586 604574
rect 478822 604338 498266 604574
rect 498502 604338 498586 604574
rect 498822 604338 518266 604574
rect 518502 604338 518586 604574
rect 518822 604338 538266 604574
rect 538502 604338 538586 604574
rect 538822 604338 558266 604574
rect 558502 604338 558586 604574
rect 558822 604338 578266 604574
rect 578502 604338 578586 604574
rect 578822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 14546 601174
rect 14782 600938 14866 601174
rect 15102 600938 34546 601174
rect 34782 600938 34866 601174
rect 35102 600938 54546 601174
rect 54782 600938 54866 601174
rect 55102 600938 74546 601174
rect 74782 600938 74866 601174
rect 75102 600938 94546 601174
rect 94782 600938 94866 601174
rect 95102 600938 114546 601174
rect 114782 600938 114866 601174
rect 115102 600938 134546 601174
rect 134782 600938 134866 601174
rect 135102 600938 154546 601174
rect 154782 600938 154866 601174
rect 155102 600938 174546 601174
rect 174782 600938 174866 601174
rect 175102 600938 194546 601174
rect 194782 600938 194866 601174
rect 195102 600938 214546 601174
rect 214782 600938 214866 601174
rect 215102 600938 234546 601174
rect 234782 600938 234866 601174
rect 235102 600938 254546 601174
rect 254782 600938 254866 601174
rect 255102 600938 274546 601174
rect 274782 600938 274866 601174
rect 275102 600938 294546 601174
rect 294782 600938 294866 601174
rect 295102 600938 314546 601174
rect 314782 600938 314866 601174
rect 315102 600938 334546 601174
rect 334782 600938 334866 601174
rect 335102 600938 354546 601174
rect 354782 600938 354866 601174
rect 355102 600938 374546 601174
rect 374782 600938 374866 601174
rect 375102 600938 394546 601174
rect 394782 600938 394866 601174
rect 395102 600938 414546 601174
rect 414782 600938 414866 601174
rect 415102 600938 434546 601174
rect 434782 600938 434866 601174
rect 435102 600938 454546 601174
rect 454782 600938 454866 601174
rect 455102 600938 474546 601174
rect 474782 600938 474866 601174
rect 475102 600938 494546 601174
rect 494782 600938 494866 601174
rect 495102 600938 514546 601174
rect 514782 600938 514866 601174
rect 515102 600938 534546 601174
rect 534782 600938 534866 601174
rect 535102 600938 554546 601174
rect 554782 600938 554866 601174
rect 555102 600938 574546 601174
rect 574782 600938 574866 601174
rect 575102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 14546 600854
rect 14782 600618 14866 600854
rect 15102 600618 34546 600854
rect 34782 600618 34866 600854
rect 35102 600618 54546 600854
rect 54782 600618 54866 600854
rect 55102 600618 74546 600854
rect 74782 600618 74866 600854
rect 75102 600618 94546 600854
rect 94782 600618 94866 600854
rect 95102 600618 114546 600854
rect 114782 600618 114866 600854
rect 115102 600618 134546 600854
rect 134782 600618 134866 600854
rect 135102 600618 154546 600854
rect 154782 600618 154866 600854
rect 155102 600618 174546 600854
rect 174782 600618 174866 600854
rect 175102 600618 194546 600854
rect 194782 600618 194866 600854
rect 195102 600618 214546 600854
rect 214782 600618 214866 600854
rect 215102 600618 234546 600854
rect 234782 600618 234866 600854
rect 235102 600618 254546 600854
rect 254782 600618 254866 600854
rect 255102 600618 274546 600854
rect 274782 600618 274866 600854
rect 275102 600618 294546 600854
rect 294782 600618 294866 600854
rect 295102 600618 314546 600854
rect 314782 600618 314866 600854
rect 315102 600618 334546 600854
rect 334782 600618 334866 600854
rect 335102 600618 354546 600854
rect 354782 600618 354866 600854
rect 355102 600618 374546 600854
rect 374782 600618 374866 600854
rect 375102 600618 394546 600854
rect 394782 600618 394866 600854
rect 395102 600618 414546 600854
rect 414782 600618 414866 600854
rect 415102 600618 434546 600854
rect 434782 600618 434866 600854
rect 435102 600618 454546 600854
rect 454782 600618 454866 600854
rect 455102 600618 474546 600854
rect 474782 600618 474866 600854
rect 475102 600618 494546 600854
rect 494782 600618 494866 600854
rect 495102 600618 514546 600854
rect 514782 600618 514866 600854
rect 515102 600618 534546 600854
rect 534782 600618 534866 600854
rect 535102 600618 554546 600854
rect 554782 600618 554866 600854
rect 555102 600618 574546 600854
rect 574782 600618 574866 600854
rect 575102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 10826 597454
rect 11062 597218 11146 597454
rect 11382 597218 30826 597454
rect 31062 597218 31146 597454
rect 31382 597218 50826 597454
rect 51062 597218 51146 597454
rect 51382 597218 70826 597454
rect 71062 597218 71146 597454
rect 71382 597218 90826 597454
rect 91062 597218 91146 597454
rect 91382 597218 110826 597454
rect 111062 597218 111146 597454
rect 111382 597218 130826 597454
rect 131062 597218 131146 597454
rect 131382 597218 150826 597454
rect 151062 597218 151146 597454
rect 151382 597218 170826 597454
rect 171062 597218 171146 597454
rect 171382 597218 190826 597454
rect 191062 597218 191146 597454
rect 191382 597218 210826 597454
rect 211062 597218 211146 597454
rect 211382 597218 230826 597454
rect 231062 597218 231146 597454
rect 231382 597218 250826 597454
rect 251062 597218 251146 597454
rect 251382 597218 270826 597454
rect 271062 597218 271146 597454
rect 271382 597218 290826 597454
rect 291062 597218 291146 597454
rect 291382 597218 310826 597454
rect 311062 597218 311146 597454
rect 311382 597218 330826 597454
rect 331062 597218 331146 597454
rect 331382 597218 350826 597454
rect 351062 597218 351146 597454
rect 351382 597218 370826 597454
rect 371062 597218 371146 597454
rect 371382 597218 390826 597454
rect 391062 597218 391146 597454
rect 391382 597218 410826 597454
rect 411062 597218 411146 597454
rect 411382 597218 430826 597454
rect 431062 597218 431146 597454
rect 431382 597218 450826 597454
rect 451062 597218 451146 597454
rect 451382 597218 470826 597454
rect 471062 597218 471146 597454
rect 471382 597218 490826 597454
rect 491062 597218 491146 597454
rect 491382 597218 510826 597454
rect 511062 597218 511146 597454
rect 511382 597218 530826 597454
rect 531062 597218 531146 597454
rect 531382 597218 550826 597454
rect 551062 597218 551146 597454
rect 551382 597218 570826 597454
rect 571062 597218 571146 597454
rect 571382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 10826 597134
rect 11062 596898 11146 597134
rect 11382 596898 30826 597134
rect 31062 596898 31146 597134
rect 31382 596898 50826 597134
rect 51062 596898 51146 597134
rect 51382 596898 70826 597134
rect 71062 596898 71146 597134
rect 71382 596898 90826 597134
rect 91062 596898 91146 597134
rect 91382 596898 110826 597134
rect 111062 596898 111146 597134
rect 111382 596898 130826 597134
rect 131062 596898 131146 597134
rect 131382 596898 150826 597134
rect 151062 596898 151146 597134
rect 151382 596898 170826 597134
rect 171062 596898 171146 597134
rect 171382 596898 190826 597134
rect 191062 596898 191146 597134
rect 191382 596898 210826 597134
rect 211062 596898 211146 597134
rect 211382 596898 230826 597134
rect 231062 596898 231146 597134
rect 231382 596898 250826 597134
rect 251062 596898 251146 597134
rect 251382 596898 270826 597134
rect 271062 596898 271146 597134
rect 271382 596898 290826 597134
rect 291062 596898 291146 597134
rect 291382 596898 310826 597134
rect 311062 596898 311146 597134
rect 311382 596898 330826 597134
rect 331062 596898 331146 597134
rect 331382 596898 350826 597134
rect 351062 596898 351146 597134
rect 351382 596898 370826 597134
rect 371062 596898 371146 597134
rect 371382 596898 390826 597134
rect 391062 596898 391146 597134
rect 391382 596898 410826 597134
rect 411062 596898 411146 597134
rect 411382 596898 430826 597134
rect 431062 596898 431146 597134
rect 431382 596898 450826 597134
rect 451062 596898 451146 597134
rect 451382 596898 470826 597134
rect 471062 596898 471146 597134
rect 471382 596898 490826 597134
rect 491062 596898 491146 597134
rect 491382 596898 510826 597134
rect 511062 596898 511146 597134
rect 511382 596898 530826 597134
rect 531062 596898 531146 597134
rect 531382 596898 550826 597134
rect 551062 596898 551146 597134
rect 551382 596898 570826 597134
rect 571062 596898 571146 597134
rect 571382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 11986 590614
rect 12222 590378 12306 590614
rect 12542 590378 31986 590614
rect 32222 590378 32306 590614
rect 32542 590378 51986 590614
rect 52222 590378 52306 590614
rect 52542 590378 71986 590614
rect 72222 590378 72306 590614
rect 72542 590378 91986 590614
rect 92222 590378 92306 590614
rect 92542 590378 111986 590614
rect 112222 590378 112306 590614
rect 112542 590378 131986 590614
rect 132222 590378 132306 590614
rect 132542 590378 151986 590614
rect 152222 590378 152306 590614
rect 152542 590378 171986 590614
rect 172222 590378 172306 590614
rect 172542 590378 191986 590614
rect 192222 590378 192306 590614
rect 192542 590378 211986 590614
rect 212222 590378 212306 590614
rect 212542 590378 231986 590614
rect 232222 590378 232306 590614
rect 232542 590378 251986 590614
rect 252222 590378 252306 590614
rect 252542 590378 271986 590614
rect 272222 590378 272306 590614
rect 272542 590378 291986 590614
rect 292222 590378 292306 590614
rect 292542 590378 311986 590614
rect 312222 590378 312306 590614
rect 312542 590378 331986 590614
rect 332222 590378 332306 590614
rect 332542 590378 351986 590614
rect 352222 590378 352306 590614
rect 352542 590378 371986 590614
rect 372222 590378 372306 590614
rect 372542 590378 391986 590614
rect 392222 590378 392306 590614
rect 392542 590378 411986 590614
rect 412222 590378 412306 590614
rect 412542 590378 431986 590614
rect 432222 590378 432306 590614
rect 432542 590378 451986 590614
rect 452222 590378 452306 590614
rect 452542 590378 471986 590614
rect 472222 590378 472306 590614
rect 472542 590378 491986 590614
rect 492222 590378 492306 590614
rect 492542 590378 511986 590614
rect 512222 590378 512306 590614
rect 512542 590378 531986 590614
rect 532222 590378 532306 590614
rect 532542 590378 551986 590614
rect 552222 590378 552306 590614
rect 552542 590378 571986 590614
rect 572222 590378 572306 590614
rect 572542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 11986 590294
rect 12222 590058 12306 590294
rect 12542 590058 31986 590294
rect 32222 590058 32306 590294
rect 32542 590058 51986 590294
rect 52222 590058 52306 590294
rect 52542 590058 71986 590294
rect 72222 590058 72306 590294
rect 72542 590058 91986 590294
rect 92222 590058 92306 590294
rect 92542 590058 111986 590294
rect 112222 590058 112306 590294
rect 112542 590058 131986 590294
rect 132222 590058 132306 590294
rect 132542 590058 151986 590294
rect 152222 590058 152306 590294
rect 152542 590058 171986 590294
rect 172222 590058 172306 590294
rect 172542 590058 191986 590294
rect 192222 590058 192306 590294
rect 192542 590058 211986 590294
rect 212222 590058 212306 590294
rect 212542 590058 231986 590294
rect 232222 590058 232306 590294
rect 232542 590058 251986 590294
rect 252222 590058 252306 590294
rect 252542 590058 271986 590294
rect 272222 590058 272306 590294
rect 272542 590058 291986 590294
rect 292222 590058 292306 590294
rect 292542 590058 311986 590294
rect 312222 590058 312306 590294
rect 312542 590058 331986 590294
rect 332222 590058 332306 590294
rect 332542 590058 351986 590294
rect 352222 590058 352306 590294
rect 352542 590058 371986 590294
rect 372222 590058 372306 590294
rect 372542 590058 391986 590294
rect 392222 590058 392306 590294
rect 392542 590058 411986 590294
rect 412222 590058 412306 590294
rect 412542 590058 431986 590294
rect 432222 590058 432306 590294
rect 432542 590058 451986 590294
rect 452222 590058 452306 590294
rect 452542 590058 471986 590294
rect 472222 590058 472306 590294
rect 472542 590058 491986 590294
rect 492222 590058 492306 590294
rect 492542 590058 511986 590294
rect 512222 590058 512306 590294
rect 512542 590058 531986 590294
rect 532222 590058 532306 590294
rect 532542 590058 551986 590294
rect 552222 590058 552306 590294
rect 552542 590058 571986 590294
rect 572222 590058 572306 590294
rect 572542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 8266 586894
rect 8502 586658 8586 586894
rect 8822 586658 28266 586894
rect 28502 586658 28586 586894
rect 28822 586658 48266 586894
rect 48502 586658 48586 586894
rect 48822 586658 68266 586894
rect 68502 586658 68586 586894
rect 68822 586658 88266 586894
rect 88502 586658 88586 586894
rect 88822 586658 108266 586894
rect 108502 586658 108586 586894
rect 108822 586658 128266 586894
rect 128502 586658 128586 586894
rect 128822 586658 148266 586894
rect 148502 586658 148586 586894
rect 148822 586658 168266 586894
rect 168502 586658 168586 586894
rect 168822 586658 188266 586894
rect 188502 586658 188586 586894
rect 188822 586658 208266 586894
rect 208502 586658 208586 586894
rect 208822 586658 228266 586894
rect 228502 586658 228586 586894
rect 228822 586658 248266 586894
rect 248502 586658 248586 586894
rect 248822 586658 268266 586894
rect 268502 586658 268586 586894
rect 268822 586658 288266 586894
rect 288502 586658 288586 586894
rect 288822 586658 308266 586894
rect 308502 586658 308586 586894
rect 308822 586658 328266 586894
rect 328502 586658 328586 586894
rect 328822 586658 348266 586894
rect 348502 586658 348586 586894
rect 348822 586658 368266 586894
rect 368502 586658 368586 586894
rect 368822 586658 388266 586894
rect 388502 586658 388586 586894
rect 388822 586658 408266 586894
rect 408502 586658 408586 586894
rect 408822 586658 428266 586894
rect 428502 586658 428586 586894
rect 428822 586658 448266 586894
rect 448502 586658 448586 586894
rect 448822 586658 468266 586894
rect 468502 586658 468586 586894
rect 468822 586658 488266 586894
rect 488502 586658 488586 586894
rect 488822 586658 508266 586894
rect 508502 586658 508586 586894
rect 508822 586658 528266 586894
rect 528502 586658 528586 586894
rect 528822 586658 548266 586894
rect 548502 586658 548586 586894
rect 548822 586658 568266 586894
rect 568502 586658 568586 586894
rect 568822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 8266 586574
rect 8502 586338 8586 586574
rect 8822 586338 28266 586574
rect 28502 586338 28586 586574
rect 28822 586338 48266 586574
rect 48502 586338 48586 586574
rect 48822 586338 68266 586574
rect 68502 586338 68586 586574
rect 68822 586338 88266 586574
rect 88502 586338 88586 586574
rect 88822 586338 108266 586574
rect 108502 586338 108586 586574
rect 108822 586338 128266 586574
rect 128502 586338 128586 586574
rect 128822 586338 148266 586574
rect 148502 586338 148586 586574
rect 148822 586338 168266 586574
rect 168502 586338 168586 586574
rect 168822 586338 188266 586574
rect 188502 586338 188586 586574
rect 188822 586338 208266 586574
rect 208502 586338 208586 586574
rect 208822 586338 228266 586574
rect 228502 586338 228586 586574
rect 228822 586338 248266 586574
rect 248502 586338 248586 586574
rect 248822 586338 268266 586574
rect 268502 586338 268586 586574
rect 268822 586338 288266 586574
rect 288502 586338 288586 586574
rect 288822 586338 308266 586574
rect 308502 586338 308586 586574
rect 308822 586338 328266 586574
rect 328502 586338 328586 586574
rect 328822 586338 348266 586574
rect 348502 586338 348586 586574
rect 348822 586338 368266 586574
rect 368502 586338 368586 586574
rect 368822 586338 388266 586574
rect 388502 586338 388586 586574
rect 388822 586338 408266 586574
rect 408502 586338 408586 586574
rect 408822 586338 428266 586574
rect 428502 586338 428586 586574
rect 428822 586338 448266 586574
rect 448502 586338 448586 586574
rect 448822 586338 468266 586574
rect 468502 586338 468586 586574
rect 468822 586338 488266 586574
rect 488502 586338 488586 586574
rect 488822 586338 508266 586574
rect 508502 586338 508586 586574
rect 508822 586338 528266 586574
rect 528502 586338 528586 586574
rect 528822 586338 548266 586574
rect 548502 586338 548586 586574
rect 548822 586338 568266 586574
rect 568502 586338 568586 586574
rect 568822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 4546 583174
rect 4782 582938 4866 583174
rect 5102 582938 24546 583174
rect 24782 582938 24866 583174
rect 25102 582938 44546 583174
rect 44782 582938 44866 583174
rect 45102 582938 64546 583174
rect 64782 582938 64866 583174
rect 65102 582938 84546 583174
rect 84782 582938 84866 583174
rect 85102 582938 104546 583174
rect 104782 582938 104866 583174
rect 105102 582938 124546 583174
rect 124782 582938 124866 583174
rect 125102 582938 144546 583174
rect 144782 582938 144866 583174
rect 145102 582938 164546 583174
rect 164782 582938 164866 583174
rect 165102 582938 184546 583174
rect 184782 582938 184866 583174
rect 185102 582938 204546 583174
rect 204782 582938 204866 583174
rect 205102 582938 224546 583174
rect 224782 582938 224866 583174
rect 225102 582938 244546 583174
rect 244782 582938 244866 583174
rect 245102 582938 264546 583174
rect 264782 582938 264866 583174
rect 265102 582938 284546 583174
rect 284782 582938 284866 583174
rect 285102 582938 304546 583174
rect 304782 582938 304866 583174
rect 305102 582938 324546 583174
rect 324782 582938 324866 583174
rect 325102 582938 344546 583174
rect 344782 582938 344866 583174
rect 345102 582938 364546 583174
rect 364782 582938 364866 583174
rect 365102 582938 384546 583174
rect 384782 582938 384866 583174
rect 385102 582938 404546 583174
rect 404782 582938 404866 583174
rect 405102 582938 424546 583174
rect 424782 582938 424866 583174
rect 425102 582938 444546 583174
rect 444782 582938 444866 583174
rect 445102 582938 464546 583174
rect 464782 582938 464866 583174
rect 465102 582938 484546 583174
rect 484782 582938 484866 583174
rect 485102 582938 504546 583174
rect 504782 582938 504866 583174
rect 505102 582938 524546 583174
rect 524782 582938 524866 583174
rect 525102 582938 544546 583174
rect 544782 582938 544866 583174
rect 545102 582938 564546 583174
rect 564782 582938 564866 583174
rect 565102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 4546 582854
rect 4782 582618 4866 582854
rect 5102 582618 24546 582854
rect 24782 582618 24866 582854
rect 25102 582618 44546 582854
rect 44782 582618 44866 582854
rect 45102 582618 64546 582854
rect 64782 582618 64866 582854
rect 65102 582618 84546 582854
rect 84782 582618 84866 582854
rect 85102 582618 104546 582854
rect 104782 582618 104866 582854
rect 105102 582618 124546 582854
rect 124782 582618 124866 582854
rect 125102 582618 144546 582854
rect 144782 582618 144866 582854
rect 145102 582618 164546 582854
rect 164782 582618 164866 582854
rect 165102 582618 184546 582854
rect 184782 582618 184866 582854
rect 185102 582618 204546 582854
rect 204782 582618 204866 582854
rect 205102 582618 224546 582854
rect 224782 582618 224866 582854
rect 225102 582618 244546 582854
rect 244782 582618 244866 582854
rect 245102 582618 264546 582854
rect 264782 582618 264866 582854
rect 265102 582618 284546 582854
rect 284782 582618 284866 582854
rect 285102 582618 304546 582854
rect 304782 582618 304866 582854
rect 305102 582618 324546 582854
rect 324782 582618 324866 582854
rect 325102 582618 344546 582854
rect 344782 582618 344866 582854
rect 345102 582618 364546 582854
rect 364782 582618 364866 582854
rect 365102 582618 384546 582854
rect 384782 582618 384866 582854
rect 385102 582618 404546 582854
rect 404782 582618 404866 582854
rect 405102 582618 424546 582854
rect 424782 582618 424866 582854
rect 425102 582618 444546 582854
rect 444782 582618 444866 582854
rect 445102 582618 464546 582854
rect 464782 582618 464866 582854
rect 465102 582618 484546 582854
rect 484782 582618 484866 582854
rect 485102 582618 504546 582854
rect 504782 582618 504866 582854
rect 505102 582618 524546 582854
rect 524782 582618 524866 582854
rect 525102 582618 544546 582854
rect 544782 582618 544866 582854
rect 545102 582618 564546 582854
rect 564782 582618 564866 582854
rect 565102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 826 579454
rect 1062 579218 1146 579454
rect 1382 579218 20826 579454
rect 21062 579218 21146 579454
rect 21382 579218 40826 579454
rect 41062 579218 41146 579454
rect 41382 579218 60826 579454
rect 61062 579218 61146 579454
rect 61382 579218 80826 579454
rect 81062 579218 81146 579454
rect 81382 579218 100826 579454
rect 101062 579218 101146 579454
rect 101382 579218 120826 579454
rect 121062 579218 121146 579454
rect 121382 579218 140826 579454
rect 141062 579218 141146 579454
rect 141382 579218 160826 579454
rect 161062 579218 161146 579454
rect 161382 579218 180826 579454
rect 181062 579218 181146 579454
rect 181382 579218 200826 579454
rect 201062 579218 201146 579454
rect 201382 579218 220826 579454
rect 221062 579218 221146 579454
rect 221382 579218 240826 579454
rect 241062 579218 241146 579454
rect 241382 579218 260826 579454
rect 261062 579218 261146 579454
rect 261382 579218 280826 579454
rect 281062 579218 281146 579454
rect 281382 579218 300826 579454
rect 301062 579218 301146 579454
rect 301382 579218 320826 579454
rect 321062 579218 321146 579454
rect 321382 579218 340826 579454
rect 341062 579218 341146 579454
rect 341382 579218 360826 579454
rect 361062 579218 361146 579454
rect 361382 579218 380826 579454
rect 381062 579218 381146 579454
rect 381382 579218 400826 579454
rect 401062 579218 401146 579454
rect 401382 579218 420826 579454
rect 421062 579218 421146 579454
rect 421382 579218 440826 579454
rect 441062 579218 441146 579454
rect 441382 579218 460826 579454
rect 461062 579218 461146 579454
rect 461382 579218 480826 579454
rect 481062 579218 481146 579454
rect 481382 579218 500826 579454
rect 501062 579218 501146 579454
rect 501382 579218 520826 579454
rect 521062 579218 521146 579454
rect 521382 579218 540826 579454
rect 541062 579218 541146 579454
rect 541382 579218 560826 579454
rect 561062 579218 561146 579454
rect 561382 579218 580826 579454
rect 581062 579218 581146 579454
rect 581382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 826 579134
rect 1062 578898 1146 579134
rect 1382 578898 20826 579134
rect 21062 578898 21146 579134
rect 21382 578898 40826 579134
rect 41062 578898 41146 579134
rect 41382 578898 60826 579134
rect 61062 578898 61146 579134
rect 61382 578898 80826 579134
rect 81062 578898 81146 579134
rect 81382 578898 100826 579134
rect 101062 578898 101146 579134
rect 101382 578898 120826 579134
rect 121062 578898 121146 579134
rect 121382 578898 140826 579134
rect 141062 578898 141146 579134
rect 141382 578898 160826 579134
rect 161062 578898 161146 579134
rect 161382 578898 180826 579134
rect 181062 578898 181146 579134
rect 181382 578898 200826 579134
rect 201062 578898 201146 579134
rect 201382 578898 220826 579134
rect 221062 578898 221146 579134
rect 221382 578898 240826 579134
rect 241062 578898 241146 579134
rect 241382 578898 260826 579134
rect 261062 578898 261146 579134
rect 261382 578898 280826 579134
rect 281062 578898 281146 579134
rect 281382 578898 300826 579134
rect 301062 578898 301146 579134
rect 301382 578898 320826 579134
rect 321062 578898 321146 579134
rect 321382 578898 340826 579134
rect 341062 578898 341146 579134
rect 341382 578898 360826 579134
rect 361062 578898 361146 579134
rect 361382 578898 380826 579134
rect 381062 578898 381146 579134
rect 381382 578898 400826 579134
rect 401062 578898 401146 579134
rect 401382 578898 420826 579134
rect 421062 578898 421146 579134
rect 421382 578898 440826 579134
rect 441062 578898 441146 579134
rect 441382 578898 460826 579134
rect 461062 578898 461146 579134
rect 461382 578898 480826 579134
rect 481062 578898 481146 579134
rect 481382 578898 500826 579134
rect 501062 578898 501146 579134
rect 501382 578898 520826 579134
rect 521062 578898 521146 579134
rect 521382 578898 540826 579134
rect 541062 578898 541146 579134
rect 541382 578898 560826 579134
rect 561062 578898 561146 579134
rect 561382 578898 580826 579134
rect 581062 578898 581146 579134
rect 581382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 21986 572614
rect 22222 572378 22306 572614
rect 22542 572378 41986 572614
rect 42222 572378 42306 572614
rect 42542 572378 61986 572614
rect 62222 572378 62306 572614
rect 62542 572378 81986 572614
rect 82222 572378 82306 572614
rect 82542 572378 101986 572614
rect 102222 572378 102306 572614
rect 102542 572378 121986 572614
rect 122222 572378 122306 572614
rect 122542 572378 141986 572614
rect 142222 572378 142306 572614
rect 142542 572378 161986 572614
rect 162222 572378 162306 572614
rect 162542 572378 181986 572614
rect 182222 572378 182306 572614
rect 182542 572378 201986 572614
rect 202222 572378 202306 572614
rect 202542 572378 221986 572614
rect 222222 572378 222306 572614
rect 222542 572378 241986 572614
rect 242222 572378 242306 572614
rect 242542 572378 261986 572614
rect 262222 572378 262306 572614
rect 262542 572378 281986 572614
rect 282222 572378 282306 572614
rect 282542 572378 301986 572614
rect 302222 572378 302306 572614
rect 302542 572378 321986 572614
rect 322222 572378 322306 572614
rect 322542 572378 341986 572614
rect 342222 572378 342306 572614
rect 342542 572378 361986 572614
rect 362222 572378 362306 572614
rect 362542 572378 381986 572614
rect 382222 572378 382306 572614
rect 382542 572378 401986 572614
rect 402222 572378 402306 572614
rect 402542 572378 421986 572614
rect 422222 572378 422306 572614
rect 422542 572378 441986 572614
rect 442222 572378 442306 572614
rect 442542 572378 461986 572614
rect 462222 572378 462306 572614
rect 462542 572378 481986 572614
rect 482222 572378 482306 572614
rect 482542 572378 501986 572614
rect 502222 572378 502306 572614
rect 502542 572378 521986 572614
rect 522222 572378 522306 572614
rect 522542 572378 541986 572614
rect 542222 572378 542306 572614
rect 542542 572378 561986 572614
rect 562222 572378 562306 572614
rect 562542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 21986 572294
rect 22222 572058 22306 572294
rect 22542 572058 41986 572294
rect 42222 572058 42306 572294
rect 42542 572058 61986 572294
rect 62222 572058 62306 572294
rect 62542 572058 81986 572294
rect 82222 572058 82306 572294
rect 82542 572058 101986 572294
rect 102222 572058 102306 572294
rect 102542 572058 121986 572294
rect 122222 572058 122306 572294
rect 122542 572058 141986 572294
rect 142222 572058 142306 572294
rect 142542 572058 161986 572294
rect 162222 572058 162306 572294
rect 162542 572058 181986 572294
rect 182222 572058 182306 572294
rect 182542 572058 201986 572294
rect 202222 572058 202306 572294
rect 202542 572058 221986 572294
rect 222222 572058 222306 572294
rect 222542 572058 241986 572294
rect 242222 572058 242306 572294
rect 242542 572058 261986 572294
rect 262222 572058 262306 572294
rect 262542 572058 281986 572294
rect 282222 572058 282306 572294
rect 282542 572058 301986 572294
rect 302222 572058 302306 572294
rect 302542 572058 321986 572294
rect 322222 572058 322306 572294
rect 322542 572058 341986 572294
rect 342222 572058 342306 572294
rect 342542 572058 361986 572294
rect 362222 572058 362306 572294
rect 362542 572058 381986 572294
rect 382222 572058 382306 572294
rect 382542 572058 401986 572294
rect 402222 572058 402306 572294
rect 402542 572058 421986 572294
rect 422222 572058 422306 572294
rect 422542 572058 441986 572294
rect 442222 572058 442306 572294
rect 442542 572058 461986 572294
rect 462222 572058 462306 572294
rect 462542 572058 481986 572294
rect 482222 572058 482306 572294
rect 482542 572058 501986 572294
rect 502222 572058 502306 572294
rect 502542 572058 521986 572294
rect 522222 572058 522306 572294
rect 522542 572058 541986 572294
rect 542222 572058 542306 572294
rect 542542 572058 561986 572294
rect 562222 572058 562306 572294
rect 562542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 18266 568894
rect 18502 568658 18586 568894
rect 18822 568658 38266 568894
rect 38502 568658 38586 568894
rect 38822 568658 58266 568894
rect 58502 568658 58586 568894
rect 58822 568658 78266 568894
rect 78502 568658 78586 568894
rect 78822 568658 98266 568894
rect 98502 568658 98586 568894
rect 98822 568658 118266 568894
rect 118502 568658 118586 568894
rect 118822 568658 138266 568894
rect 138502 568658 138586 568894
rect 138822 568658 158266 568894
rect 158502 568658 158586 568894
rect 158822 568658 178266 568894
rect 178502 568658 178586 568894
rect 178822 568658 198266 568894
rect 198502 568658 198586 568894
rect 198822 568658 218266 568894
rect 218502 568658 218586 568894
rect 218822 568658 238266 568894
rect 238502 568658 238586 568894
rect 238822 568658 258266 568894
rect 258502 568658 258586 568894
rect 258822 568658 278266 568894
rect 278502 568658 278586 568894
rect 278822 568658 298266 568894
rect 298502 568658 298586 568894
rect 298822 568658 318266 568894
rect 318502 568658 318586 568894
rect 318822 568658 338266 568894
rect 338502 568658 338586 568894
rect 338822 568658 358266 568894
rect 358502 568658 358586 568894
rect 358822 568658 378266 568894
rect 378502 568658 378586 568894
rect 378822 568658 398266 568894
rect 398502 568658 398586 568894
rect 398822 568658 418266 568894
rect 418502 568658 418586 568894
rect 418822 568658 438266 568894
rect 438502 568658 438586 568894
rect 438822 568658 458266 568894
rect 458502 568658 458586 568894
rect 458822 568658 478266 568894
rect 478502 568658 478586 568894
rect 478822 568658 498266 568894
rect 498502 568658 498586 568894
rect 498822 568658 518266 568894
rect 518502 568658 518586 568894
rect 518822 568658 538266 568894
rect 538502 568658 538586 568894
rect 538822 568658 558266 568894
rect 558502 568658 558586 568894
rect 558822 568658 578266 568894
rect 578502 568658 578586 568894
rect 578822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 18266 568574
rect 18502 568338 18586 568574
rect 18822 568338 38266 568574
rect 38502 568338 38586 568574
rect 38822 568338 58266 568574
rect 58502 568338 58586 568574
rect 58822 568338 78266 568574
rect 78502 568338 78586 568574
rect 78822 568338 98266 568574
rect 98502 568338 98586 568574
rect 98822 568338 118266 568574
rect 118502 568338 118586 568574
rect 118822 568338 138266 568574
rect 138502 568338 138586 568574
rect 138822 568338 158266 568574
rect 158502 568338 158586 568574
rect 158822 568338 178266 568574
rect 178502 568338 178586 568574
rect 178822 568338 198266 568574
rect 198502 568338 198586 568574
rect 198822 568338 218266 568574
rect 218502 568338 218586 568574
rect 218822 568338 238266 568574
rect 238502 568338 238586 568574
rect 238822 568338 258266 568574
rect 258502 568338 258586 568574
rect 258822 568338 278266 568574
rect 278502 568338 278586 568574
rect 278822 568338 298266 568574
rect 298502 568338 298586 568574
rect 298822 568338 318266 568574
rect 318502 568338 318586 568574
rect 318822 568338 338266 568574
rect 338502 568338 338586 568574
rect 338822 568338 358266 568574
rect 358502 568338 358586 568574
rect 358822 568338 378266 568574
rect 378502 568338 378586 568574
rect 378822 568338 398266 568574
rect 398502 568338 398586 568574
rect 398822 568338 418266 568574
rect 418502 568338 418586 568574
rect 418822 568338 438266 568574
rect 438502 568338 438586 568574
rect 438822 568338 458266 568574
rect 458502 568338 458586 568574
rect 458822 568338 478266 568574
rect 478502 568338 478586 568574
rect 478822 568338 498266 568574
rect 498502 568338 498586 568574
rect 498822 568338 518266 568574
rect 518502 568338 518586 568574
rect 518822 568338 538266 568574
rect 538502 568338 538586 568574
rect 538822 568338 558266 568574
rect 558502 568338 558586 568574
rect 558822 568338 578266 568574
rect 578502 568338 578586 568574
rect 578822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 14546 565174
rect 14782 564938 14866 565174
rect 15102 564938 34546 565174
rect 34782 564938 34866 565174
rect 35102 564938 54546 565174
rect 54782 564938 54866 565174
rect 55102 564938 74546 565174
rect 74782 564938 74866 565174
rect 75102 564938 94546 565174
rect 94782 564938 94866 565174
rect 95102 564938 114546 565174
rect 114782 564938 114866 565174
rect 115102 564938 134546 565174
rect 134782 564938 134866 565174
rect 135102 564938 154546 565174
rect 154782 564938 154866 565174
rect 155102 564938 174546 565174
rect 174782 564938 174866 565174
rect 175102 564938 194546 565174
rect 194782 564938 194866 565174
rect 195102 564938 214546 565174
rect 214782 564938 214866 565174
rect 215102 564938 234546 565174
rect 234782 564938 234866 565174
rect 235102 564938 254546 565174
rect 254782 564938 254866 565174
rect 255102 564938 274546 565174
rect 274782 564938 274866 565174
rect 275102 564938 294546 565174
rect 294782 564938 294866 565174
rect 295102 564938 314546 565174
rect 314782 564938 314866 565174
rect 315102 564938 334546 565174
rect 334782 564938 334866 565174
rect 335102 564938 354546 565174
rect 354782 564938 354866 565174
rect 355102 564938 374546 565174
rect 374782 564938 374866 565174
rect 375102 564938 394546 565174
rect 394782 564938 394866 565174
rect 395102 564938 414546 565174
rect 414782 564938 414866 565174
rect 415102 564938 434546 565174
rect 434782 564938 434866 565174
rect 435102 564938 454546 565174
rect 454782 564938 454866 565174
rect 455102 564938 474546 565174
rect 474782 564938 474866 565174
rect 475102 564938 494546 565174
rect 494782 564938 494866 565174
rect 495102 564938 514546 565174
rect 514782 564938 514866 565174
rect 515102 564938 534546 565174
rect 534782 564938 534866 565174
rect 535102 564938 554546 565174
rect 554782 564938 554866 565174
rect 555102 564938 574546 565174
rect 574782 564938 574866 565174
rect 575102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 14546 564854
rect 14782 564618 14866 564854
rect 15102 564618 34546 564854
rect 34782 564618 34866 564854
rect 35102 564618 54546 564854
rect 54782 564618 54866 564854
rect 55102 564618 74546 564854
rect 74782 564618 74866 564854
rect 75102 564618 94546 564854
rect 94782 564618 94866 564854
rect 95102 564618 114546 564854
rect 114782 564618 114866 564854
rect 115102 564618 134546 564854
rect 134782 564618 134866 564854
rect 135102 564618 154546 564854
rect 154782 564618 154866 564854
rect 155102 564618 174546 564854
rect 174782 564618 174866 564854
rect 175102 564618 194546 564854
rect 194782 564618 194866 564854
rect 195102 564618 214546 564854
rect 214782 564618 214866 564854
rect 215102 564618 234546 564854
rect 234782 564618 234866 564854
rect 235102 564618 254546 564854
rect 254782 564618 254866 564854
rect 255102 564618 274546 564854
rect 274782 564618 274866 564854
rect 275102 564618 294546 564854
rect 294782 564618 294866 564854
rect 295102 564618 314546 564854
rect 314782 564618 314866 564854
rect 315102 564618 334546 564854
rect 334782 564618 334866 564854
rect 335102 564618 354546 564854
rect 354782 564618 354866 564854
rect 355102 564618 374546 564854
rect 374782 564618 374866 564854
rect 375102 564618 394546 564854
rect 394782 564618 394866 564854
rect 395102 564618 414546 564854
rect 414782 564618 414866 564854
rect 415102 564618 434546 564854
rect 434782 564618 434866 564854
rect 435102 564618 454546 564854
rect 454782 564618 454866 564854
rect 455102 564618 474546 564854
rect 474782 564618 474866 564854
rect 475102 564618 494546 564854
rect 494782 564618 494866 564854
rect 495102 564618 514546 564854
rect 514782 564618 514866 564854
rect 515102 564618 534546 564854
rect 534782 564618 534866 564854
rect 535102 564618 554546 564854
rect 554782 564618 554866 564854
rect 555102 564618 574546 564854
rect 574782 564618 574866 564854
rect 575102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 10826 561454
rect 11062 561218 11146 561454
rect 11382 561218 30826 561454
rect 31062 561218 31146 561454
rect 31382 561218 50826 561454
rect 51062 561218 51146 561454
rect 51382 561218 70826 561454
rect 71062 561218 71146 561454
rect 71382 561218 90826 561454
rect 91062 561218 91146 561454
rect 91382 561218 110826 561454
rect 111062 561218 111146 561454
rect 111382 561218 130826 561454
rect 131062 561218 131146 561454
rect 131382 561218 150826 561454
rect 151062 561218 151146 561454
rect 151382 561218 170826 561454
rect 171062 561218 171146 561454
rect 171382 561218 190826 561454
rect 191062 561218 191146 561454
rect 191382 561218 210826 561454
rect 211062 561218 211146 561454
rect 211382 561218 230826 561454
rect 231062 561218 231146 561454
rect 231382 561218 250826 561454
rect 251062 561218 251146 561454
rect 251382 561218 270826 561454
rect 271062 561218 271146 561454
rect 271382 561218 290826 561454
rect 291062 561218 291146 561454
rect 291382 561218 310826 561454
rect 311062 561218 311146 561454
rect 311382 561218 330826 561454
rect 331062 561218 331146 561454
rect 331382 561218 350826 561454
rect 351062 561218 351146 561454
rect 351382 561218 370826 561454
rect 371062 561218 371146 561454
rect 371382 561218 390826 561454
rect 391062 561218 391146 561454
rect 391382 561218 410826 561454
rect 411062 561218 411146 561454
rect 411382 561218 430826 561454
rect 431062 561218 431146 561454
rect 431382 561218 450826 561454
rect 451062 561218 451146 561454
rect 451382 561218 470826 561454
rect 471062 561218 471146 561454
rect 471382 561218 490826 561454
rect 491062 561218 491146 561454
rect 491382 561218 510826 561454
rect 511062 561218 511146 561454
rect 511382 561218 530826 561454
rect 531062 561218 531146 561454
rect 531382 561218 550826 561454
rect 551062 561218 551146 561454
rect 551382 561218 570826 561454
rect 571062 561218 571146 561454
rect 571382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 10826 561134
rect 11062 560898 11146 561134
rect 11382 560898 30826 561134
rect 31062 560898 31146 561134
rect 31382 560898 50826 561134
rect 51062 560898 51146 561134
rect 51382 560898 70826 561134
rect 71062 560898 71146 561134
rect 71382 560898 90826 561134
rect 91062 560898 91146 561134
rect 91382 560898 110826 561134
rect 111062 560898 111146 561134
rect 111382 560898 130826 561134
rect 131062 560898 131146 561134
rect 131382 560898 150826 561134
rect 151062 560898 151146 561134
rect 151382 560898 170826 561134
rect 171062 560898 171146 561134
rect 171382 560898 190826 561134
rect 191062 560898 191146 561134
rect 191382 560898 210826 561134
rect 211062 560898 211146 561134
rect 211382 560898 230826 561134
rect 231062 560898 231146 561134
rect 231382 560898 250826 561134
rect 251062 560898 251146 561134
rect 251382 560898 270826 561134
rect 271062 560898 271146 561134
rect 271382 560898 290826 561134
rect 291062 560898 291146 561134
rect 291382 560898 310826 561134
rect 311062 560898 311146 561134
rect 311382 560898 330826 561134
rect 331062 560898 331146 561134
rect 331382 560898 350826 561134
rect 351062 560898 351146 561134
rect 351382 560898 370826 561134
rect 371062 560898 371146 561134
rect 371382 560898 390826 561134
rect 391062 560898 391146 561134
rect 391382 560898 410826 561134
rect 411062 560898 411146 561134
rect 411382 560898 430826 561134
rect 431062 560898 431146 561134
rect 431382 560898 450826 561134
rect 451062 560898 451146 561134
rect 451382 560898 470826 561134
rect 471062 560898 471146 561134
rect 471382 560898 490826 561134
rect 491062 560898 491146 561134
rect 491382 560898 510826 561134
rect 511062 560898 511146 561134
rect 511382 560898 530826 561134
rect 531062 560898 531146 561134
rect 531382 560898 550826 561134
rect 551062 560898 551146 561134
rect 551382 560898 570826 561134
rect 571062 560898 571146 561134
rect 571382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 11986 554614
rect 12222 554378 12306 554614
rect 12542 554378 31986 554614
rect 32222 554378 32306 554614
rect 32542 554378 51986 554614
rect 52222 554378 52306 554614
rect 52542 554378 71986 554614
rect 72222 554378 72306 554614
rect 72542 554378 91986 554614
rect 92222 554378 92306 554614
rect 92542 554378 111986 554614
rect 112222 554378 112306 554614
rect 112542 554378 131986 554614
rect 132222 554378 132306 554614
rect 132542 554378 151986 554614
rect 152222 554378 152306 554614
rect 152542 554378 171986 554614
rect 172222 554378 172306 554614
rect 172542 554378 191986 554614
rect 192222 554378 192306 554614
rect 192542 554378 211986 554614
rect 212222 554378 212306 554614
rect 212542 554378 231986 554614
rect 232222 554378 232306 554614
rect 232542 554378 251986 554614
rect 252222 554378 252306 554614
rect 252542 554378 271986 554614
rect 272222 554378 272306 554614
rect 272542 554378 291986 554614
rect 292222 554378 292306 554614
rect 292542 554378 311986 554614
rect 312222 554378 312306 554614
rect 312542 554378 331986 554614
rect 332222 554378 332306 554614
rect 332542 554378 351986 554614
rect 352222 554378 352306 554614
rect 352542 554378 371986 554614
rect 372222 554378 372306 554614
rect 372542 554378 391986 554614
rect 392222 554378 392306 554614
rect 392542 554378 411986 554614
rect 412222 554378 412306 554614
rect 412542 554378 431986 554614
rect 432222 554378 432306 554614
rect 432542 554378 451986 554614
rect 452222 554378 452306 554614
rect 452542 554378 471986 554614
rect 472222 554378 472306 554614
rect 472542 554378 491986 554614
rect 492222 554378 492306 554614
rect 492542 554378 511986 554614
rect 512222 554378 512306 554614
rect 512542 554378 531986 554614
rect 532222 554378 532306 554614
rect 532542 554378 551986 554614
rect 552222 554378 552306 554614
rect 552542 554378 571986 554614
rect 572222 554378 572306 554614
rect 572542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 11986 554294
rect 12222 554058 12306 554294
rect 12542 554058 31986 554294
rect 32222 554058 32306 554294
rect 32542 554058 51986 554294
rect 52222 554058 52306 554294
rect 52542 554058 71986 554294
rect 72222 554058 72306 554294
rect 72542 554058 91986 554294
rect 92222 554058 92306 554294
rect 92542 554058 111986 554294
rect 112222 554058 112306 554294
rect 112542 554058 131986 554294
rect 132222 554058 132306 554294
rect 132542 554058 151986 554294
rect 152222 554058 152306 554294
rect 152542 554058 171986 554294
rect 172222 554058 172306 554294
rect 172542 554058 191986 554294
rect 192222 554058 192306 554294
rect 192542 554058 211986 554294
rect 212222 554058 212306 554294
rect 212542 554058 231986 554294
rect 232222 554058 232306 554294
rect 232542 554058 251986 554294
rect 252222 554058 252306 554294
rect 252542 554058 271986 554294
rect 272222 554058 272306 554294
rect 272542 554058 291986 554294
rect 292222 554058 292306 554294
rect 292542 554058 311986 554294
rect 312222 554058 312306 554294
rect 312542 554058 331986 554294
rect 332222 554058 332306 554294
rect 332542 554058 351986 554294
rect 352222 554058 352306 554294
rect 352542 554058 371986 554294
rect 372222 554058 372306 554294
rect 372542 554058 391986 554294
rect 392222 554058 392306 554294
rect 392542 554058 411986 554294
rect 412222 554058 412306 554294
rect 412542 554058 431986 554294
rect 432222 554058 432306 554294
rect 432542 554058 451986 554294
rect 452222 554058 452306 554294
rect 452542 554058 471986 554294
rect 472222 554058 472306 554294
rect 472542 554058 491986 554294
rect 492222 554058 492306 554294
rect 492542 554058 511986 554294
rect 512222 554058 512306 554294
rect 512542 554058 531986 554294
rect 532222 554058 532306 554294
rect 532542 554058 551986 554294
rect 552222 554058 552306 554294
rect 552542 554058 571986 554294
rect 572222 554058 572306 554294
rect 572542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 8266 550894
rect 8502 550658 8586 550894
rect 8822 550658 28266 550894
rect 28502 550658 28586 550894
rect 28822 550658 48266 550894
rect 48502 550658 48586 550894
rect 48822 550658 68266 550894
rect 68502 550658 68586 550894
rect 68822 550658 88266 550894
rect 88502 550658 88586 550894
rect 88822 550658 108266 550894
rect 108502 550658 108586 550894
rect 108822 550658 128266 550894
rect 128502 550658 128586 550894
rect 128822 550658 148266 550894
rect 148502 550658 148586 550894
rect 148822 550658 168266 550894
rect 168502 550658 168586 550894
rect 168822 550658 188266 550894
rect 188502 550658 188586 550894
rect 188822 550658 208266 550894
rect 208502 550658 208586 550894
rect 208822 550658 228266 550894
rect 228502 550658 228586 550894
rect 228822 550658 248266 550894
rect 248502 550658 248586 550894
rect 248822 550658 268266 550894
rect 268502 550658 268586 550894
rect 268822 550658 288266 550894
rect 288502 550658 288586 550894
rect 288822 550658 308266 550894
rect 308502 550658 308586 550894
rect 308822 550658 328266 550894
rect 328502 550658 328586 550894
rect 328822 550658 348266 550894
rect 348502 550658 348586 550894
rect 348822 550658 368266 550894
rect 368502 550658 368586 550894
rect 368822 550658 388266 550894
rect 388502 550658 388586 550894
rect 388822 550658 408266 550894
rect 408502 550658 408586 550894
rect 408822 550658 428266 550894
rect 428502 550658 428586 550894
rect 428822 550658 448266 550894
rect 448502 550658 448586 550894
rect 448822 550658 468266 550894
rect 468502 550658 468586 550894
rect 468822 550658 488266 550894
rect 488502 550658 488586 550894
rect 488822 550658 508266 550894
rect 508502 550658 508586 550894
rect 508822 550658 528266 550894
rect 528502 550658 528586 550894
rect 528822 550658 548266 550894
rect 548502 550658 548586 550894
rect 548822 550658 568266 550894
rect 568502 550658 568586 550894
rect 568822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 8266 550574
rect 8502 550338 8586 550574
rect 8822 550338 28266 550574
rect 28502 550338 28586 550574
rect 28822 550338 48266 550574
rect 48502 550338 48586 550574
rect 48822 550338 68266 550574
rect 68502 550338 68586 550574
rect 68822 550338 88266 550574
rect 88502 550338 88586 550574
rect 88822 550338 108266 550574
rect 108502 550338 108586 550574
rect 108822 550338 128266 550574
rect 128502 550338 128586 550574
rect 128822 550338 148266 550574
rect 148502 550338 148586 550574
rect 148822 550338 168266 550574
rect 168502 550338 168586 550574
rect 168822 550338 188266 550574
rect 188502 550338 188586 550574
rect 188822 550338 208266 550574
rect 208502 550338 208586 550574
rect 208822 550338 228266 550574
rect 228502 550338 228586 550574
rect 228822 550338 248266 550574
rect 248502 550338 248586 550574
rect 248822 550338 268266 550574
rect 268502 550338 268586 550574
rect 268822 550338 288266 550574
rect 288502 550338 288586 550574
rect 288822 550338 308266 550574
rect 308502 550338 308586 550574
rect 308822 550338 328266 550574
rect 328502 550338 328586 550574
rect 328822 550338 348266 550574
rect 348502 550338 348586 550574
rect 348822 550338 368266 550574
rect 368502 550338 368586 550574
rect 368822 550338 388266 550574
rect 388502 550338 388586 550574
rect 388822 550338 408266 550574
rect 408502 550338 408586 550574
rect 408822 550338 428266 550574
rect 428502 550338 428586 550574
rect 428822 550338 448266 550574
rect 448502 550338 448586 550574
rect 448822 550338 468266 550574
rect 468502 550338 468586 550574
rect 468822 550338 488266 550574
rect 488502 550338 488586 550574
rect 488822 550338 508266 550574
rect 508502 550338 508586 550574
rect 508822 550338 528266 550574
rect 528502 550338 528586 550574
rect 528822 550338 548266 550574
rect 548502 550338 548586 550574
rect 548822 550338 568266 550574
rect 568502 550338 568586 550574
rect 568822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 4546 547174
rect 4782 546938 4866 547174
rect 5102 546938 24546 547174
rect 24782 546938 24866 547174
rect 25102 546938 44546 547174
rect 44782 546938 44866 547174
rect 45102 546938 64546 547174
rect 64782 546938 64866 547174
rect 65102 546938 84546 547174
rect 84782 546938 84866 547174
rect 85102 546938 104546 547174
rect 104782 546938 104866 547174
rect 105102 546938 124546 547174
rect 124782 546938 124866 547174
rect 125102 546938 144546 547174
rect 144782 546938 144866 547174
rect 145102 546938 164546 547174
rect 164782 546938 164866 547174
rect 165102 546938 184546 547174
rect 184782 546938 184866 547174
rect 185102 546938 204546 547174
rect 204782 546938 204866 547174
rect 205102 546938 224546 547174
rect 224782 546938 224866 547174
rect 225102 546938 244546 547174
rect 244782 546938 244866 547174
rect 245102 546938 264546 547174
rect 264782 546938 264866 547174
rect 265102 546938 284546 547174
rect 284782 546938 284866 547174
rect 285102 546938 304546 547174
rect 304782 546938 304866 547174
rect 305102 546938 324546 547174
rect 324782 546938 324866 547174
rect 325102 546938 344546 547174
rect 344782 546938 344866 547174
rect 345102 546938 364546 547174
rect 364782 546938 364866 547174
rect 365102 546938 384546 547174
rect 384782 546938 384866 547174
rect 385102 546938 404546 547174
rect 404782 546938 404866 547174
rect 405102 546938 424546 547174
rect 424782 546938 424866 547174
rect 425102 546938 444546 547174
rect 444782 546938 444866 547174
rect 445102 546938 464546 547174
rect 464782 546938 464866 547174
rect 465102 546938 484546 547174
rect 484782 546938 484866 547174
rect 485102 546938 504546 547174
rect 504782 546938 504866 547174
rect 505102 546938 524546 547174
rect 524782 546938 524866 547174
rect 525102 546938 544546 547174
rect 544782 546938 544866 547174
rect 545102 546938 564546 547174
rect 564782 546938 564866 547174
rect 565102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 4546 546854
rect 4782 546618 4866 546854
rect 5102 546618 24546 546854
rect 24782 546618 24866 546854
rect 25102 546618 44546 546854
rect 44782 546618 44866 546854
rect 45102 546618 64546 546854
rect 64782 546618 64866 546854
rect 65102 546618 84546 546854
rect 84782 546618 84866 546854
rect 85102 546618 104546 546854
rect 104782 546618 104866 546854
rect 105102 546618 124546 546854
rect 124782 546618 124866 546854
rect 125102 546618 144546 546854
rect 144782 546618 144866 546854
rect 145102 546618 164546 546854
rect 164782 546618 164866 546854
rect 165102 546618 184546 546854
rect 184782 546618 184866 546854
rect 185102 546618 204546 546854
rect 204782 546618 204866 546854
rect 205102 546618 224546 546854
rect 224782 546618 224866 546854
rect 225102 546618 244546 546854
rect 244782 546618 244866 546854
rect 245102 546618 264546 546854
rect 264782 546618 264866 546854
rect 265102 546618 284546 546854
rect 284782 546618 284866 546854
rect 285102 546618 304546 546854
rect 304782 546618 304866 546854
rect 305102 546618 324546 546854
rect 324782 546618 324866 546854
rect 325102 546618 344546 546854
rect 344782 546618 344866 546854
rect 345102 546618 364546 546854
rect 364782 546618 364866 546854
rect 365102 546618 384546 546854
rect 384782 546618 384866 546854
rect 385102 546618 404546 546854
rect 404782 546618 404866 546854
rect 405102 546618 424546 546854
rect 424782 546618 424866 546854
rect 425102 546618 444546 546854
rect 444782 546618 444866 546854
rect 445102 546618 464546 546854
rect 464782 546618 464866 546854
rect 465102 546618 484546 546854
rect 484782 546618 484866 546854
rect 485102 546618 504546 546854
rect 504782 546618 504866 546854
rect 505102 546618 524546 546854
rect 524782 546618 524866 546854
rect 525102 546618 544546 546854
rect 544782 546618 544866 546854
rect 545102 546618 564546 546854
rect 564782 546618 564866 546854
rect 565102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 826 543454
rect 1062 543218 1146 543454
rect 1382 543218 20826 543454
rect 21062 543218 21146 543454
rect 21382 543218 40826 543454
rect 41062 543218 41146 543454
rect 41382 543218 60826 543454
rect 61062 543218 61146 543454
rect 61382 543218 80826 543454
rect 81062 543218 81146 543454
rect 81382 543218 100826 543454
rect 101062 543218 101146 543454
rect 101382 543218 120826 543454
rect 121062 543218 121146 543454
rect 121382 543218 140826 543454
rect 141062 543218 141146 543454
rect 141382 543218 160826 543454
rect 161062 543218 161146 543454
rect 161382 543218 180826 543454
rect 181062 543218 181146 543454
rect 181382 543218 200826 543454
rect 201062 543218 201146 543454
rect 201382 543218 220826 543454
rect 221062 543218 221146 543454
rect 221382 543218 240826 543454
rect 241062 543218 241146 543454
rect 241382 543218 260826 543454
rect 261062 543218 261146 543454
rect 261382 543218 280826 543454
rect 281062 543218 281146 543454
rect 281382 543218 300826 543454
rect 301062 543218 301146 543454
rect 301382 543218 320826 543454
rect 321062 543218 321146 543454
rect 321382 543218 340826 543454
rect 341062 543218 341146 543454
rect 341382 543218 360826 543454
rect 361062 543218 361146 543454
rect 361382 543218 380826 543454
rect 381062 543218 381146 543454
rect 381382 543218 400826 543454
rect 401062 543218 401146 543454
rect 401382 543218 420826 543454
rect 421062 543218 421146 543454
rect 421382 543218 440826 543454
rect 441062 543218 441146 543454
rect 441382 543218 460826 543454
rect 461062 543218 461146 543454
rect 461382 543218 480826 543454
rect 481062 543218 481146 543454
rect 481382 543218 500826 543454
rect 501062 543218 501146 543454
rect 501382 543218 520826 543454
rect 521062 543218 521146 543454
rect 521382 543218 540826 543454
rect 541062 543218 541146 543454
rect 541382 543218 560826 543454
rect 561062 543218 561146 543454
rect 561382 543218 580826 543454
rect 581062 543218 581146 543454
rect 581382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 826 543134
rect 1062 542898 1146 543134
rect 1382 542898 20826 543134
rect 21062 542898 21146 543134
rect 21382 542898 40826 543134
rect 41062 542898 41146 543134
rect 41382 542898 60826 543134
rect 61062 542898 61146 543134
rect 61382 542898 80826 543134
rect 81062 542898 81146 543134
rect 81382 542898 100826 543134
rect 101062 542898 101146 543134
rect 101382 542898 120826 543134
rect 121062 542898 121146 543134
rect 121382 542898 140826 543134
rect 141062 542898 141146 543134
rect 141382 542898 160826 543134
rect 161062 542898 161146 543134
rect 161382 542898 180826 543134
rect 181062 542898 181146 543134
rect 181382 542898 200826 543134
rect 201062 542898 201146 543134
rect 201382 542898 220826 543134
rect 221062 542898 221146 543134
rect 221382 542898 240826 543134
rect 241062 542898 241146 543134
rect 241382 542898 260826 543134
rect 261062 542898 261146 543134
rect 261382 542898 280826 543134
rect 281062 542898 281146 543134
rect 281382 542898 300826 543134
rect 301062 542898 301146 543134
rect 301382 542898 320826 543134
rect 321062 542898 321146 543134
rect 321382 542898 340826 543134
rect 341062 542898 341146 543134
rect 341382 542898 360826 543134
rect 361062 542898 361146 543134
rect 361382 542898 380826 543134
rect 381062 542898 381146 543134
rect 381382 542898 400826 543134
rect 401062 542898 401146 543134
rect 401382 542898 420826 543134
rect 421062 542898 421146 543134
rect 421382 542898 440826 543134
rect 441062 542898 441146 543134
rect 441382 542898 460826 543134
rect 461062 542898 461146 543134
rect 461382 542898 480826 543134
rect 481062 542898 481146 543134
rect 481382 542898 500826 543134
rect 501062 542898 501146 543134
rect 501382 542898 520826 543134
rect 521062 542898 521146 543134
rect 521382 542898 540826 543134
rect 541062 542898 541146 543134
rect 541382 542898 560826 543134
rect 561062 542898 561146 543134
rect 561382 542898 580826 543134
rect 581062 542898 581146 543134
rect 581382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 21986 536614
rect 22222 536378 22306 536614
rect 22542 536378 41986 536614
rect 42222 536378 42306 536614
rect 42542 536378 61986 536614
rect 62222 536378 62306 536614
rect 62542 536378 81986 536614
rect 82222 536378 82306 536614
rect 82542 536378 101986 536614
rect 102222 536378 102306 536614
rect 102542 536378 121986 536614
rect 122222 536378 122306 536614
rect 122542 536378 141986 536614
rect 142222 536378 142306 536614
rect 142542 536378 161986 536614
rect 162222 536378 162306 536614
rect 162542 536378 181986 536614
rect 182222 536378 182306 536614
rect 182542 536378 201986 536614
rect 202222 536378 202306 536614
rect 202542 536378 221986 536614
rect 222222 536378 222306 536614
rect 222542 536378 241986 536614
rect 242222 536378 242306 536614
rect 242542 536378 261986 536614
rect 262222 536378 262306 536614
rect 262542 536378 281986 536614
rect 282222 536378 282306 536614
rect 282542 536378 301986 536614
rect 302222 536378 302306 536614
rect 302542 536378 321986 536614
rect 322222 536378 322306 536614
rect 322542 536378 341986 536614
rect 342222 536378 342306 536614
rect 342542 536378 361986 536614
rect 362222 536378 362306 536614
rect 362542 536378 381986 536614
rect 382222 536378 382306 536614
rect 382542 536378 401986 536614
rect 402222 536378 402306 536614
rect 402542 536378 421986 536614
rect 422222 536378 422306 536614
rect 422542 536378 441986 536614
rect 442222 536378 442306 536614
rect 442542 536378 461986 536614
rect 462222 536378 462306 536614
rect 462542 536378 481986 536614
rect 482222 536378 482306 536614
rect 482542 536378 501986 536614
rect 502222 536378 502306 536614
rect 502542 536378 521986 536614
rect 522222 536378 522306 536614
rect 522542 536378 541986 536614
rect 542222 536378 542306 536614
rect 542542 536378 561986 536614
rect 562222 536378 562306 536614
rect 562542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 21986 536294
rect 22222 536058 22306 536294
rect 22542 536058 41986 536294
rect 42222 536058 42306 536294
rect 42542 536058 61986 536294
rect 62222 536058 62306 536294
rect 62542 536058 81986 536294
rect 82222 536058 82306 536294
rect 82542 536058 101986 536294
rect 102222 536058 102306 536294
rect 102542 536058 121986 536294
rect 122222 536058 122306 536294
rect 122542 536058 141986 536294
rect 142222 536058 142306 536294
rect 142542 536058 161986 536294
rect 162222 536058 162306 536294
rect 162542 536058 181986 536294
rect 182222 536058 182306 536294
rect 182542 536058 201986 536294
rect 202222 536058 202306 536294
rect 202542 536058 221986 536294
rect 222222 536058 222306 536294
rect 222542 536058 241986 536294
rect 242222 536058 242306 536294
rect 242542 536058 261986 536294
rect 262222 536058 262306 536294
rect 262542 536058 281986 536294
rect 282222 536058 282306 536294
rect 282542 536058 301986 536294
rect 302222 536058 302306 536294
rect 302542 536058 321986 536294
rect 322222 536058 322306 536294
rect 322542 536058 341986 536294
rect 342222 536058 342306 536294
rect 342542 536058 361986 536294
rect 362222 536058 362306 536294
rect 362542 536058 381986 536294
rect 382222 536058 382306 536294
rect 382542 536058 401986 536294
rect 402222 536058 402306 536294
rect 402542 536058 421986 536294
rect 422222 536058 422306 536294
rect 422542 536058 441986 536294
rect 442222 536058 442306 536294
rect 442542 536058 461986 536294
rect 462222 536058 462306 536294
rect 462542 536058 481986 536294
rect 482222 536058 482306 536294
rect 482542 536058 501986 536294
rect 502222 536058 502306 536294
rect 502542 536058 521986 536294
rect 522222 536058 522306 536294
rect 522542 536058 541986 536294
rect 542222 536058 542306 536294
rect 542542 536058 561986 536294
rect 562222 536058 562306 536294
rect 562542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 18266 532894
rect 18502 532658 18586 532894
rect 18822 532658 38266 532894
rect 38502 532658 38586 532894
rect 38822 532658 58266 532894
rect 58502 532658 58586 532894
rect 58822 532658 78266 532894
rect 78502 532658 78586 532894
rect 78822 532658 98266 532894
rect 98502 532658 98586 532894
rect 98822 532658 118266 532894
rect 118502 532658 118586 532894
rect 118822 532658 138266 532894
rect 138502 532658 138586 532894
rect 138822 532658 158266 532894
rect 158502 532658 158586 532894
rect 158822 532658 178266 532894
rect 178502 532658 178586 532894
rect 178822 532658 198266 532894
rect 198502 532658 198586 532894
rect 198822 532658 218266 532894
rect 218502 532658 218586 532894
rect 218822 532658 238266 532894
rect 238502 532658 238586 532894
rect 238822 532658 258266 532894
rect 258502 532658 258586 532894
rect 258822 532658 278266 532894
rect 278502 532658 278586 532894
rect 278822 532658 298266 532894
rect 298502 532658 298586 532894
rect 298822 532658 318266 532894
rect 318502 532658 318586 532894
rect 318822 532658 338266 532894
rect 338502 532658 338586 532894
rect 338822 532658 358266 532894
rect 358502 532658 358586 532894
rect 358822 532658 378266 532894
rect 378502 532658 378586 532894
rect 378822 532658 398266 532894
rect 398502 532658 398586 532894
rect 398822 532658 418266 532894
rect 418502 532658 418586 532894
rect 418822 532658 438266 532894
rect 438502 532658 438586 532894
rect 438822 532658 458266 532894
rect 458502 532658 458586 532894
rect 458822 532658 478266 532894
rect 478502 532658 478586 532894
rect 478822 532658 498266 532894
rect 498502 532658 498586 532894
rect 498822 532658 518266 532894
rect 518502 532658 518586 532894
rect 518822 532658 538266 532894
rect 538502 532658 538586 532894
rect 538822 532658 558266 532894
rect 558502 532658 558586 532894
rect 558822 532658 578266 532894
rect 578502 532658 578586 532894
rect 578822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 18266 532574
rect 18502 532338 18586 532574
rect 18822 532338 38266 532574
rect 38502 532338 38586 532574
rect 38822 532338 58266 532574
rect 58502 532338 58586 532574
rect 58822 532338 78266 532574
rect 78502 532338 78586 532574
rect 78822 532338 98266 532574
rect 98502 532338 98586 532574
rect 98822 532338 118266 532574
rect 118502 532338 118586 532574
rect 118822 532338 138266 532574
rect 138502 532338 138586 532574
rect 138822 532338 158266 532574
rect 158502 532338 158586 532574
rect 158822 532338 178266 532574
rect 178502 532338 178586 532574
rect 178822 532338 198266 532574
rect 198502 532338 198586 532574
rect 198822 532338 218266 532574
rect 218502 532338 218586 532574
rect 218822 532338 238266 532574
rect 238502 532338 238586 532574
rect 238822 532338 258266 532574
rect 258502 532338 258586 532574
rect 258822 532338 278266 532574
rect 278502 532338 278586 532574
rect 278822 532338 298266 532574
rect 298502 532338 298586 532574
rect 298822 532338 318266 532574
rect 318502 532338 318586 532574
rect 318822 532338 338266 532574
rect 338502 532338 338586 532574
rect 338822 532338 358266 532574
rect 358502 532338 358586 532574
rect 358822 532338 378266 532574
rect 378502 532338 378586 532574
rect 378822 532338 398266 532574
rect 398502 532338 398586 532574
rect 398822 532338 418266 532574
rect 418502 532338 418586 532574
rect 418822 532338 438266 532574
rect 438502 532338 438586 532574
rect 438822 532338 458266 532574
rect 458502 532338 458586 532574
rect 458822 532338 478266 532574
rect 478502 532338 478586 532574
rect 478822 532338 498266 532574
rect 498502 532338 498586 532574
rect 498822 532338 518266 532574
rect 518502 532338 518586 532574
rect 518822 532338 538266 532574
rect 538502 532338 538586 532574
rect 538822 532338 558266 532574
rect 558502 532338 558586 532574
rect 558822 532338 578266 532574
rect 578502 532338 578586 532574
rect 578822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 14546 529174
rect 14782 528938 14866 529174
rect 15102 528938 34546 529174
rect 34782 528938 34866 529174
rect 35102 528938 54546 529174
rect 54782 528938 54866 529174
rect 55102 528938 74546 529174
rect 74782 528938 74866 529174
rect 75102 528938 94546 529174
rect 94782 528938 94866 529174
rect 95102 528938 114546 529174
rect 114782 528938 114866 529174
rect 115102 528938 134546 529174
rect 134782 528938 134866 529174
rect 135102 528938 154546 529174
rect 154782 528938 154866 529174
rect 155102 528938 174546 529174
rect 174782 528938 174866 529174
rect 175102 528938 194546 529174
rect 194782 528938 194866 529174
rect 195102 528938 214546 529174
rect 214782 528938 214866 529174
rect 215102 528938 234546 529174
rect 234782 528938 234866 529174
rect 235102 528938 254546 529174
rect 254782 528938 254866 529174
rect 255102 528938 274546 529174
rect 274782 528938 274866 529174
rect 275102 528938 294546 529174
rect 294782 528938 294866 529174
rect 295102 528938 314546 529174
rect 314782 528938 314866 529174
rect 315102 528938 334546 529174
rect 334782 528938 334866 529174
rect 335102 528938 354546 529174
rect 354782 528938 354866 529174
rect 355102 528938 374546 529174
rect 374782 528938 374866 529174
rect 375102 528938 394546 529174
rect 394782 528938 394866 529174
rect 395102 528938 414546 529174
rect 414782 528938 414866 529174
rect 415102 528938 434546 529174
rect 434782 528938 434866 529174
rect 435102 528938 454546 529174
rect 454782 528938 454866 529174
rect 455102 528938 474546 529174
rect 474782 528938 474866 529174
rect 475102 528938 494546 529174
rect 494782 528938 494866 529174
rect 495102 528938 514546 529174
rect 514782 528938 514866 529174
rect 515102 528938 534546 529174
rect 534782 528938 534866 529174
rect 535102 528938 554546 529174
rect 554782 528938 554866 529174
rect 555102 528938 574546 529174
rect 574782 528938 574866 529174
rect 575102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 14546 528854
rect 14782 528618 14866 528854
rect 15102 528618 34546 528854
rect 34782 528618 34866 528854
rect 35102 528618 54546 528854
rect 54782 528618 54866 528854
rect 55102 528618 74546 528854
rect 74782 528618 74866 528854
rect 75102 528618 94546 528854
rect 94782 528618 94866 528854
rect 95102 528618 114546 528854
rect 114782 528618 114866 528854
rect 115102 528618 134546 528854
rect 134782 528618 134866 528854
rect 135102 528618 154546 528854
rect 154782 528618 154866 528854
rect 155102 528618 174546 528854
rect 174782 528618 174866 528854
rect 175102 528618 194546 528854
rect 194782 528618 194866 528854
rect 195102 528618 214546 528854
rect 214782 528618 214866 528854
rect 215102 528618 234546 528854
rect 234782 528618 234866 528854
rect 235102 528618 254546 528854
rect 254782 528618 254866 528854
rect 255102 528618 274546 528854
rect 274782 528618 274866 528854
rect 275102 528618 294546 528854
rect 294782 528618 294866 528854
rect 295102 528618 314546 528854
rect 314782 528618 314866 528854
rect 315102 528618 334546 528854
rect 334782 528618 334866 528854
rect 335102 528618 354546 528854
rect 354782 528618 354866 528854
rect 355102 528618 374546 528854
rect 374782 528618 374866 528854
rect 375102 528618 394546 528854
rect 394782 528618 394866 528854
rect 395102 528618 414546 528854
rect 414782 528618 414866 528854
rect 415102 528618 434546 528854
rect 434782 528618 434866 528854
rect 435102 528618 454546 528854
rect 454782 528618 454866 528854
rect 455102 528618 474546 528854
rect 474782 528618 474866 528854
rect 475102 528618 494546 528854
rect 494782 528618 494866 528854
rect 495102 528618 514546 528854
rect 514782 528618 514866 528854
rect 515102 528618 534546 528854
rect 534782 528618 534866 528854
rect 535102 528618 554546 528854
rect 554782 528618 554866 528854
rect 555102 528618 574546 528854
rect 574782 528618 574866 528854
rect 575102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 10826 525454
rect 11062 525218 11146 525454
rect 11382 525218 30826 525454
rect 31062 525218 31146 525454
rect 31382 525218 50826 525454
rect 51062 525218 51146 525454
rect 51382 525218 70826 525454
rect 71062 525218 71146 525454
rect 71382 525218 90826 525454
rect 91062 525218 91146 525454
rect 91382 525218 110826 525454
rect 111062 525218 111146 525454
rect 111382 525218 130826 525454
rect 131062 525218 131146 525454
rect 131382 525218 150826 525454
rect 151062 525218 151146 525454
rect 151382 525218 170826 525454
rect 171062 525218 171146 525454
rect 171382 525218 190826 525454
rect 191062 525218 191146 525454
rect 191382 525218 210826 525454
rect 211062 525218 211146 525454
rect 211382 525218 230826 525454
rect 231062 525218 231146 525454
rect 231382 525218 250826 525454
rect 251062 525218 251146 525454
rect 251382 525218 270826 525454
rect 271062 525218 271146 525454
rect 271382 525218 290826 525454
rect 291062 525218 291146 525454
rect 291382 525218 310826 525454
rect 311062 525218 311146 525454
rect 311382 525218 330826 525454
rect 331062 525218 331146 525454
rect 331382 525218 350826 525454
rect 351062 525218 351146 525454
rect 351382 525218 370826 525454
rect 371062 525218 371146 525454
rect 371382 525218 390826 525454
rect 391062 525218 391146 525454
rect 391382 525218 410826 525454
rect 411062 525218 411146 525454
rect 411382 525218 430826 525454
rect 431062 525218 431146 525454
rect 431382 525218 450826 525454
rect 451062 525218 451146 525454
rect 451382 525218 470826 525454
rect 471062 525218 471146 525454
rect 471382 525218 490826 525454
rect 491062 525218 491146 525454
rect 491382 525218 510826 525454
rect 511062 525218 511146 525454
rect 511382 525218 530826 525454
rect 531062 525218 531146 525454
rect 531382 525218 550826 525454
rect 551062 525218 551146 525454
rect 551382 525218 570826 525454
rect 571062 525218 571146 525454
rect 571382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 10826 525134
rect 11062 524898 11146 525134
rect 11382 524898 30826 525134
rect 31062 524898 31146 525134
rect 31382 524898 50826 525134
rect 51062 524898 51146 525134
rect 51382 524898 70826 525134
rect 71062 524898 71146 525134
rect 71382 524898 90826 525134
rect 91062 524898 91146 525134
rect 91382 524898 110826 525134
rect 111062 524898 111146 525134
rect 111382 524898 130826 525134
rect 131062 524898 131146 525134
rect 131382 524898 150826 525134
rect 151062 524898 151146 525134
rect 151382 524898 170826 525134
rect 171062 524898 171146 525134
rect 171382 524898 190826 525134
rect 191062 524898 191146 525134
rect 191382 524898 210826 525134
rect 211062 524898 211146 525134
rect 211382 524898 230826 525134
rect 231062 524898 231146 525134
rect 231382 524898 250826 525134
rect 251062 524898 251146 525134
rect 251382 524898 270826 525134
rect 271062 524898 271146 525134
rect 271382 524898 290826 525134
rect 291062 524898 291146 525134
rect 291382 524898 310826 525134
rect 311062 524898 311146 525134
rect 311382 524898 330826 525134
rect 331062 524898 331146 525134
rect 331382 524898 350826 525134
rect 351062 524898 351146 525134
rect 351382 524898 370826 525134
rect 371062 524898 371146 525134
rect 371382 524898 390826 525134
rect 391062 524898 391146 525134
rect 391382 524898 410826 525134
rect 411062 524898 411146 525134
rect 411382 524898 430826 525134
rect 431062 524898 431146 525134
rect 431382 524898 450826 525134
rect 451062 524898 451146 525134
rect 451382 524898 470826 525134
rect 471062 524898 471146 525134
rect 471382 524898 490826 525134
rect 491062 524898 491146 525134
rect 491382 524898 510826 525134
rect 511062 524898 511146 525134
rect 511382 524898 530826 525134
rect 531062 524898 531146 525134
rect 531382 524898 550826 525134
rect 551062 524898 551146 525134
rect 551382 524898 570826 525134
rect 571062 524898 571146 525134
rect 571382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 11986 518614
rect 12222 518378 12306 518614
rect 12542 518378 31986 518614
rect 32222 518378 32306 518614
rect 32542 518378 51986 518614
rect 52222 518378 52306 518614
rect 52542 518378 71986 518614
rect 72222 518378 72306 518614
rect 72542 518378 91986 518614
rect 92222 518378 92306 518614
rect 92542 518378 111986 518614
rect 112222 518378 112306 518614
rect 112542 518378 131986 518614
rect 132222 518378 132306 518614
rect 132542 518378 151986 518614
rect 152222 518378 152306 518614
rect 152542 518378 171986 518614
rect 172222 518378 172306 518614
rect 172542 518378 191986 518614
rect 192222 518378 192306 518614
rect 192542 518378 211986 518614
rect 212222 518378 212306 518614
rect 212542 518378 231986 518614
rect 232222 518378 232306 518614
rect 232542 518378 251986 518614
rect 252222 518378 252306 518614
rect 252542 518378 271986 518614
rect 272222 518378 272306 518614
rect 272542 518378 291986 518614
rect 292222 518378 292306 518614
rect 292542 518378 311986 518614
rect 312222 518378 312306 518614
rect 312542 518378 331986 518614
rect 332222 518378 332306 518614
rect 332542 518378 351986 518614
rect 352222 518378 352306 518614
rect 352542 518378 371986 518614
rect 372222 518378 372306 518614
rect 372542 518378 391986 518614
rect 392222 518378 392306 518614
rect 392542 518378 411986 518614
rect 412222 518378 412306 518614
rect 412542 518378 431986 518614
rect 432222 518378 432306 518614
rect 432542 518378 451986 518614
rect 452222 518378 452306 518614
rect 452542 518378 471986 518614
rect 472222 518378 472306 518614
rect 472542 518378 491986 518614
rect 492222 518378 492306 518614
rect 492542 518378 511986 518614
rect 512222 518378 512306 518614
rect 512542 518378 531986 518614
rect 532222 518378 532306 518614
rect 532542 518378 551986 518614
rect 552222 518378 552306 518614
rect 552542 518378 571986 518614
rect 572222 518378 572306 518614
rect 572542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 11986 518294
rect 12222 518058 12306 518294
rect 12542 518058 31986 518294
rect 32222 518058 32306 518294
rect 32542 518058 51986 518294
rect 52222 518058 52306 518294
rect 52542 518058 71986 518294
rect 72222 518058 72306 518294
rect 72542 518058 91986 518294
rect 92222 518058 92306 518294
rect 92542 518058 111986 518294
rect 112222 518058 112306 518294
rect 112542 518058 131986 518294
rect 132222 518058 132306 518294
rect 132542 518058 151986 518294
rect 152222 518058 152306 518294
rect 152542 518058 171986 518294
rect 172222 518058 172306 518294
rect 172542 518058 191986 518294
rect 192222 518058 192306 518294
rect 192542 518058 211986 518294
rect 212222 518058 212306 518294
rect 212542 518058 231986 518294
rect 232222 518058 232306 518294
rect 232542 518058 251986 518294
rect 252222 518058 252306 518294
rect 252542 518058 271986 518294
rect 272222 518058 272306 518294
rect 272542 518058 291986 518294
rect 292222 518058 292306 518294
rect 292542 518058 311986 518294
rect 312222 518058 312306 518294
rect 312542 518058 331986 518294
rect 332222 518058 332306 518294
rect 332542 518058 351986 518294
rect 352222 518058 352306 518294
rect 352542 518058 371986 518294
rect 372222 518058 372306 518294
rect 372542 518058 391986 518294
rect 392222 518058 392306 518294
rect 392542 518058 411986 518294
rect 412222 518058 412306 518294
rect 412542 518058 431986 518294
rect 432222 518058 432306 518294
rect 432542 518058 451986 518294
rect 452222 518058 452306 518294
rect 452542 518058 471986 518294
rect 472222 518058 472306 518294
rect 472542 518058 491986 518294
rect 492222 518058 492306 518294
rect 492542 518058 511986 518294
rect 512222 518058 512306 518294
rect 512542 518058 531986 518294
rect 532222 518058 532306 518294
rect 532542 518058 551986 518294
rect 552222 518058 552306 518294
rect 552542 518058 571986 518294
rect 572222 518058 572306 518294
rect 572542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 8266 514894
rect 8502 514658 8586 514894
rect 8822 514658 28266 514894
rect 28502 514658 28586 514894
rect 28822 514658 48266 514894
rect 48502 514658 48586 514894
rect 48822 514658 68266 514894
rect 68502 514658 68586 514894
rect 68822 514658 88266 514894
rect 88502 514658 88586 514894
rect 88822 514658 108266 514894
rect 108502 514658 108586 514894
rect 108822 514658 128266 514894
rect 128502 514658 128586 514894
rect 128822 514658 148266 514894
rect 148502 514658 148586 514894
rect 148822 514658 168266 514894
rect 168502 514658 168586 514894
rect 168822 514658 188266 514894
rect 188502 514658 188586 514894
rect 188822 514658 208266 514894
rect 208502 514658 208586 514894
rect 208822 514658 228266 514894
rect 228502 514658 228586 514894
rect 228822 514658 248266 514894
rect 248502 514658 248586 514894
rect 248822 514658 268266 514894
rect 268502 514658 268586 514894
rect 268822 514658 288266 514894
rect 288502 514658 288586 514894
rect 288822 514658 308266 514894
rect 308502 514658 308586 514894
rect 308822 514658 328266 514894
rect 328502 514658 328586 514894
rect 328822 514658 348266 514894
rect 348502 514658 348586 514894
rect 348822 514658 368266 514894
rect 368502 514658 368586 514894
rect 368822 514658 388266 514894
rect 388502 514658 388586 514894
rect 388822 514658 408266 514894
rect 408502 514658 408586 514894
rect 408822 514658 428266 514894
rect 428502 514658 428586 514894
rect 428822 514658 448266 514894
rect 448502 514658 448586 514894
rect 448822 514658 468266 514894
rect 468502 514658 468586 514894
rect 468822 514658 488266 514894
rect 488502 514658 488586 514894
rect 488822 514658 508266 514894
rect 508502 514658 508586 514894
rect 508822 514658 528266 514894
rect 528502 514658 528586 514894
rect 528822 514658 548266 514894
rect 548502 514658 548586 514894
rect 548822 514658 568266 514894
rect 568502 514658 568586 514894
rect 568822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 8266 514574
rect 8502 514338 8586 514574
rect 8822 514338 28266 514574
rect 28502 514338 28586 514574
rect 28822 514338 48266 514574
rect 48502 514338 48586 514574
rect 48822 514338 68266 514574
rect 68502 514338 68586 514574
rect 68822 514338 88266 514574
rect 88502 514338 88586 514574
rect 88822 514338 108266 514574
rect 108502 514338 108586 514574
rect 108822 514338 128266 514574
rect 128502 514338 128586 514574
rect 128822 514338 148266 514574
rect 148502 514338 148586 514574
rect 148822 514338 168266 514574
rect 168502 514338 168586 514574
rect 168822 514338 188266 514574
rect 188502 514338 188586 514574
rect 188822 514338 208266 514574
rect 208502 514338 208586 514574
rect 208822 514338 228266 514574
rect 228502 514338 228586 514574
rect 228822 514338 248266 514574
rect 248502 514338 248586 514574
rect 248822 514338 268266 514574
rect 268502 514338 268586 514574
rect 268822 514338 288266 514574
rect 288502 514338 288586 514574
rect 288822 514338 308266 514574
rect 308502 514338 308586 514574
rect 308822 514338 328266 514574
rect 328502 514338 328586 514574
rect 328822 514338 348266 514574
rect 348502 514338 348586 514574
rect 348822 514338 368266 514574
rect 368502 514338 368586 514574
rect 368822 514338 388266 514574
rect 388502 514338 388586 514574
rect 388822 514338 408266 514574
rect 408502 514338 408586 514574
rect 408822 514338 428266 514574
rect 428502 514338 428586 514574
rect 428822 514338 448266 514574
rect 448502 514338 448586 514574
rect 448822 514338 468266 514574
rect 468502 514338 468586 514574
rect 468822 514338 488266 514574
rect 488502 514338 488586 514574
rect 488822 514338 508266 514574
rect 508502 514338 508586 514574
rect 508822 514338 528266 514574
rect 528502 514338 528586 514574
rect 528822 514338 548266 514574
rect 548502 514338 548586 514574
rect 548822 514338 568266 514574
rect 568502 514338 568586 514574
rect 568822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 4546 511174
rect 4782 510938 4866 511174
rect 5102 510938 24546 511174
rect 24782 510938 24866 511174
rect 25102 510938 44546 511174
rect 44782 510938 44866 511174
rect 45102 510938 64546 511174
rect 64782 510938 64866 511174
rect 65102 510938 84546 511174
rect 84782 510938 84866 511174
rect 85102 510938 104546 511174
rect 104782 510938 104866 511174
rect 105102 510938 124546 511174
rect 124782 510938 124866 511174
rect 125102 510938 144546 511174
rect 144782 510938 144866 511174
rect 145102 510938 164546 511174
rect 164782 510938 164866 511174
rect 165102 510938 184546 511174
rect 184782 510938 184866 511174
rect 185102 510938 204546 511174
rect 204782 510938 204866 511174
rect 205102 510938 224546 511174
rect 224782 510938 224866 511174
rect 225102 510938 244546 511174
rect 244782 510938 244866 511174
rect 245102 510938 264546 511174
rect 264782 510938 264866 511174
rect 265102 510938 284546 511174
rect 284782 510938 284866 511174
rect 285102 510938 304546 511174
rect 304782 510938 304866 511174
rect 305102 510938 324546 511174
rect 324782 510938 324866 511174
rect 325102 510938 344546 511174
rect 344782 510938 344866 511174
rect 345102 510938 364546 511174
rect 364782 510938 364866 511174
rect 365102 510938 384546 511174
rect 384782 510938 384866 511174
rect 385102 510938 404546 511174
rect 404782 510938 404866 511174
rect 405102 510938 424546 511174
rect 424782 510938 424866 511174
rect 425102 510938 444546 511174
rect 444782 510938 444866 511174
rect 445102 510938 464546 511174
rect 464782 510938 464866 511174
rect 465102 510938 484546 511174
rect 484782 510938 484866 511174
rect 485102 510938 504546 511174
rect 504782 510938 504866 511174
rect 505102 510938 524546 511174
rect 524782 510938 524866 511174
rect 525102 510938 544546 511174
rect 544782 510938 544866 511174
rect 545102 510938 564546 511174
rect 564782 510938 564866 511174
rect 565102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 4546 510854
rect 4782 510618 4866 510854
rect 5102 510618 24546 510854
rect 24782 510618 24866 510854
rect 25102 510618 44546 510854
rect 44782 510618 44866 510854
rect 45102 510618 64546 510854
rect 64782 510618 64866 510854
rect 65102 510618 84546 510854
rect 84782 510618 84866 510854
rect 85102 510618 104546 510854
rect 104782 510618 104866 510854
rect 105102 510618 124546 510854
rect 124782 510618 124866 510854
rect 125102 510618 144546 510854
rect 144782 510618 144866 510854
rect 145102 510618 164546 510854
rect 164782 510618 164866 510854
rect 165102 510618 184546 510854
rect 184782 510618 184866 510854
rect 185102 510618 204546 510854
rect 204782 510618 204866 510854
rect 205102 510618 224546 510854
rect 224782 510618 224866 510854
rect 225102 510618 244546 510854
rect 244782 510618 244866 510854
rect 245102 510618 264546 510854
rect 264782 510618 264866 510854
rect 265102 510618 284546 510854
rect 284782 510618 284866 510854
rect 285102 510618 304546 510854
rect 304782 510618 304866 510854
rect 305102 510618 324546 510854
rect 324782 510618 324866 510854
rect 325102 510618 344546 510854
rect 344782 510618 344866 510854
rect 345102 510618 364546 510854
rect 364782 510618 364866 510854
rect 365102 510618 384546 510854
rect 384782 510618 384866 510854
rect 385102 510618 404546 510854
rect 404782 510618 404866 510854
rect 405102 510618 424546 510854
rect 424782 510618 424866 510854
rect 425102 510618 444546 510854
rect 444782 510618 444866 510854
rect 445102 510618 464546 510854
rect 464782 510618 464866 510854
rect 465102 510618 484546 510854
rect 484782 510618 484866 510854
rect 485102 510618 504546 510854
rect 504782 510618 504866 510854
rect 505102 510618 524546 510854
rect 524782 510618 524866 510854
rect 525102 510618 544546 510854
rect 544782 510618 544866 510854
rect 545102 510618 564546 510854
rect 564782 510618 564866 510854
rect 565102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 826 507454
rect 1062 507218 1146 507454
rect 1382 507218 20826 507454
rect 21062 507218 21146 507454
rect 21382 507218 40826 507454
rect 41062 507218 41146 507454
rect 41382 507218 60826 507454
rect 61062 507218 61146 507454
rect 61382 507218 80826 507454
rect 81062 507218 81146 507454
rect 81382 507218 100826 507454
rect 101062 507218 101146 507454
rect 101382 507218 120826 507454
rect 121062 507218 121146 507454
rect 121382 507218 140826 507454
rect 141062 507218 141146 507454
rect 141382 507218 160826 507454
rect 161062 507218 161146 507454
rect 161382 507218 180826 507454
rect 181062 507218 181146 507454
rect 181382 507218 200826 507454
rect 201062 507218 201146 507454
rect 201382 507218 220826 507454
rect 221062 507218 221146 507454
rect 221382 507218 240826 507454
rect 241062 507218 241146 507454
rect 241382 507218 260826 507454
rect 261062 507218 261146 507454
rect 261382 507218 280826 507454
rect 281062 507218 281146 507454
rect 281382 507218 300826 507454
rect 301062 507218 301146 507454
rect 301382 507218 320826 507454
rect 321062 507218 321146 507454
rect 321382 507218 340826 507454
rect 341062 507218 341146 507454
rect 341382 507218 360826 507454
rect 361062 507218 361146 507454
rect 361382 507218 380826 507454
rect 381062 507218 381146 507454
rect 381382 507218 400826 507454
rect 401062 507218 401146 507454
rect 401382 507218 420826 507454
rect 421062 507218 421146 507454
rect 421382 507218 440826 507454
rect 441062 507218 441146 507454
rect 441382 507218 460826 507454
rect 461062 507218 461146 507454
rect 461382 507218 480826 507454
rect 481062 507218 481146 507454
rect 481382 507218 500826 507454
rect 501062 507218 501146 507454
rect 501382 507218 520826 507454
rect 521062 507218 521146 507454
rect 521382 507218 540826 507454
rect 541062 507218 541146 507454
rect 541382 507218 560826 507454
rect 561062 507218 561146 507454
rect 561382 507218 580826 507454
rect 581062 507218 581146 507454
rect 581382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 826 507134
rect 1062 506898 1146 507134
rect 1382 506898 20826 507134
rect 21062 506898 21146 507134
rect 21382 506898 40826 507134
rect 41062 506898 41146 507134
rect 41382 506898 60826 507134
rect 61062 506898 61146 507134
rect 61382 506898 80826 507134
rect 81062 506898 81146 507134
rect 81382 506898 100826 507134
rect 101062 506898 101146 507134
rect 101382 506898 120826 507134
rect 121062 506898 121146 507134
rect 121382 506898 140826 507134
rect 141062 506898 141146 507134
rect 141382 506898 160826 507134
rect 161062 506898 161146 507134
rect 161382 506898 180826 507134
rect 181062 506898 181146 507134
rect 181382 506898 200826 507134
rect 201062 506898 201146 507134
rect 201382 506898 220826 507134
rect 221062 506898 221146 507134
rect 221382 506898 240826 507134
rect 241062 506898 241146 507134
rect 241382 506898 260826 507134
rect 261062 506898 261146 507134
rect 261382 506898 280826 507134
rect 281062 506898 281146 507134
rect 281382 506898 300826 507134
rect 301062 506898 301146 507134
rect 301382 506898 320826 507134
rect 321062 506898 321146 507134
rect 321382 506898 340826 507134
rect 341062 506898 341146 507134
rect 341382 506898 360826 507134
rect 361062 506898 361146 507134
rect 361382 506898 380826 507134
rect 381062 506898 381146 507134
rect 381382 506898 400826 507134
rect 401062 506898 401146 507134
rect 401382 506898 420826 507134
rect 421062 506898 421146 507134
rect 421382 506898 440826 507134
rect 441062 506898 441146 507134
rect 441382 506898 460826 507134
rect 461062 506898 461146 507134
rect 461382 506898 480826 507134
rect 481062 506898 481146 507134
rect 481382 506898 500826 507134
rect 501062 506898 501146 507134
rect 501382 506898 520826 507134
rect 521062 506898 521146 507134
rect 521382 506898 540826 507134
rect 541062 506898 541146 507134
rect 541382 506898 560826 507134
rect 561062 506898 561146 507134
rect 561382 506898 580826 507134
rect 581062 506898 581146 507134
rect 581382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 21986 500614
rect 22222 500378 22306 500614
rect 22542 500378 41986 500614
rect 42222 500378 42306 500614
rect 42542 500378 61986 500614
rect 62222 500378 62306 500614
rect 62542 500378 81986 500614
rect 82222 500378 82306 500614
rect 82542 500378 101986 500614
rect 102222 500378 102306 500614
rect 102542 500378 121986 500614
rect 122222 500378 122306 500614
rect 122542 500378 141986 500614
rect 142222 500378 142306 500614
rect 142542 500378 161986 500614
rect 162222 500378 162306 500614
rect 162542 500378 181986 500614
rect 182222 500378 182306 500614
rect 182542 500378 201986 500614
rect 202222 500378 202306 500614
rect 202542 500378 221986 500614
rect 222222 500378 222306 500614
rect 222542 500378 241986 500614
rect 242222 500378 242306 500614
rect 242542 500378 261986 500614
rect 262222 500378 262306 500614
rect 262542 500378 281986 500614
rect 282222 500378 282306 500614
rect 282542 500378 301986 500614
rect 302222 500378 302306 500614
rect 302542 500378 321986 500614
rect 322222 500378 322306 500614
rect 322542 500378 341986 500614
rect 342222 500378 342306 500614
rect 342542 500378 361986 500614
rect 362222 500378 362306 500614
rect 362542 500378 381986 500614
rect 382222 500378 382306 500614
rect 382542 500378 401986 500614
rect 402222 500378 402306 500614
rect 402542 500378 421986 500614
rect 422222 500378 422306 500614
rect 422542 500378 441986 500614
rect 442222 500378 442306 500614
rect 442542 500378 461986 500614
rect 462222 500378 462306 500614
rect 462542 500378 481986 500614
rect 482222 500378 482306 500614
rect 482542 500378 501986 500614
rect 502222 500378 502306 500614
rect 502542 500378 521986 500614
rect 522222 500378 522306 500614
rect 522542 500378 541986 500614
rect 542222 500378 542306 500614
rect 542542 500378 561986 500614
rect 562222 500378 562306 500614
rect 562542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 21986 500294
rect 22222 500058 22306 500294
rect 22542 500058 41986 500294
rect 42222 500058 42306 500294
rect 42542 500058 61986 500294
rect 62222 500058 62306 500294
rect 62542 500058 81986 500294
rect 82222 500058 82306 500294
rect 82542 500058 101986 500294
rect 102222 500058 102306 500294
rect 102542 500058 121986 500294
rect 122222 500058 122306 500294
rect 122542 500058 141986 500294
rect 142222 500058 142306 500294
rect 142542 500058 161986 500294
rect 162222 500058 162306 500294
rect 162542 500058 181986 500294
rect 182222 500058 182306 500294
rect 182542 500058 201986 500294
rect 202222 500058 202306 500294
rect 202542 500058 221986 500294
rect 222222 500058 222306 500294
rect 222542 500058 241986 500294
rect 242222 500058 242306 500294
rect 242542 500058 261986 500294
rect 262222 500058 262306 500294
rect 262542 500058 281986 500294
rect 282222 500058 282306 500294
rect 282542 500058 301986 500294
rect 302222 500058 302306 500294
rect 302542 500058 321986 500294
rect 322222 500058 322306 500294
rect 322542 500058 341986 500294
rect 342222 500058 342306 500294
rect 342542 500058 361986 500294
rect 362222 500058 362306 500294
rect 362542 500058 381986 500294
rect 382222 500058 382306 500294
rect 382542 500058 401986 500294
rect 402222 500058 402306 500294
rect 402542 500058 421986 500294
rect 422222 500058 422306 500294
rect 422542 500058 441986 500294
rect 442222 500058 442306 500294
rect 442542 500058 461986 500294
rect 462222 500058 462306 500294
rect 462542 500058 481986 500294
rect 482222 500058 482306 500294
rect 482542 500058 501986 500294
rect 502222 500058 502306 500294
rect 502542 500058 521986 500294
rect 522222 500058 522306 500294
rect 522542 500058 541986 500294
rect 542222 500058 542306 500294
rect 542542 500058 561986 500294
rect 562222 500058 562306 500294
rect 562542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 18266 496894
rect 18502 496658 18586 496894
rect 18822 496658 38266 496894
rect 38502 496658 38586 496894
rect 38822 496658 58266 496894
rect 58502 496658 58586 496894
rect 58822 496658 78266 496894
rect 78502 496658 78586 496894
rect 78822 496658 98266 496894
rect 98502 496658 98586 496894
rect 98822 496658 118266 496894
rect 118502 496658 118586 496894
rect 118822 496658 138266 496894
rect 138502 496658 138586 496894
rect 138822 496658 158266 496894
rect 158502 496658 158586 496894
rect 158822 496658 178266 496894
rect 178502 496658 178586 496894
rect 178822 496658 198266 496894
rect 198502 496658 198586 496894
rect 198822 496658 218266 496894
rect 218502 496658 218586 496894
rect 218822 496658 238266 496894
rect 238502 496658 238586 496894
rect 238822 496658 258266 496894
rect 258502 496658 258586 496894
rect 258822 496658 278266 496894
rect 278502 496658 278586 496894
rect 278822 496658 298266 496894
rect 298502 496658 298586 496894
rect 298822 496658 318266 496894
rect 318502 496658 318586 496894
rect 318822 496658 338266 496894
rect 338502 496658 338586 496894
rect 338822 496658 358266 496894
rect 358502 496658 358586 496894
rect 358822 496658 378266 496894
rect 378502 496658 378586 496894
rect 378822 496658 398266 496894
rect 398502 496658 398586 496894
rect 398822 496658 418266 496894
rect 418502 496658 418586 496894
rect 418822 496658 438266 496894
rect 438502 496658 438586 496894
rect 438822 496658 458266 496894
rect 458502 496658 458586 496894
rect 458822 496658 478266 496894
rect 478502 496658 478586 496894
rect 478822 496658 498266 496894
rect 498502 496658 498586 496894
rect 498822 496658 518266 496894
rect 518502 496658 518586 496894
rect 518822 496658 538266 496894
rect 538502 496658 538586 496894
rect 538822 496658 558266 496894
rect 558502 496658 558586 496894
rect 558822 496658 578266 496894
rect 578502 496658 578586 496894
rect 578822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 18266 496574
rect 18502 496338 18586 496574
rect 18822 496338 38266 496574
rect 38502 496338 38586 496574
rect 38822 496338 58266 496574
rect 58502 496338 58586 496574
rect 58822 496338 78266 496574
rect 78502 496338 78586 496574
rect 78822 496338 98266 496574
rect 98502 496338 98586 496574
rect 98822 496338 118266 496574
rect 118502 496338 118586 496574
rect 118822 496338 138266 496574
rect 138502 496338 138586 496574
rect 138822 496338 158266 496574
rect 158502 496338 158586 496574
rect 158822 496338 178266 496574
rect 178502 496338 178586 496574
rect 178822 496338 198266 496574
rect 198502 496338 198586 496574
rect 198822 496338 218266 496574
rect 218502 496338 218586 496574
rect 218822 496338 238266 496574
rect 238502 496338 238586 496574
rect 238822 496338 258266 496574
rect 258502 496338 258586 496574
rect 258822 496338 278266 496574
rect 278502 496338 278586 496574
rect 278822 496338 298266 496574
rect 298502 496338 298586 496574
rect 298822 496338 318266 496574
rect 318502 496338 318586 496574
rect 318822 496338 338266 496574
rect 338502 496338 338586 496574
rect 338822 496338 358266 496574
rect 358502 496338 358586 496574
rect 358822 496338 378266 496574
rect 378502 496338 378586 496574
rect 378822 496338 398266 496574
rect 398502 496338 398586 496574
rect 398822 496338 418266 496574
rect 418502 496338 418586 496574
rect 418822 496338 438266 496574
rect 438502 496338 438586 496574
rect 438822 496338 458266 496574
rect 458502 496338 458586 496574
rect 458822 496338 478266 496574
rect 478502 496338 478586 496574
rect 478822 496338 498266 496574
rect 498502 496338 498586 496574
rect 498822 496338 518266 496574
rect 518502 496338 518586 496574
rect 518822 496338 538266 496574
rect 538502 496338 538586 496574
rect 538822 496338 558266 496574
rect 558502 496338 558586 496574
rect 558822 496338 578266 496574
rect 578502 496338 578586 496574
rect 578822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 14546 493174
rect 14782 492938 14866 493174
rect 15102 492938 34546 493174
rect 34782 492938 34866 493174
rect 35102 492938 54546 493174
rect 54782 492938 54866 493174
rect 55102 492938 74546 493174
rect 74782 492938 74866 493174
rect 75102 492938 94546 493174
rect 94782 492938 94866 493174
rect 95102 492938 114546 493174
rect 114782 492938 114866 493174
rect 115102 492938 134546 493174
rect 134782 492938 134866 493174
rect 135102 492938 154546 493174
rect 154782 492938 154866 493174
rect 155102 492938 174546 493174
rect 174782 492938 174866 493174
rect 175102 492938 194546 493174
rect 194782 492938 194866 493174
rect 195102 492938 214546 493174
rect 214782 492938 214866 493174
rect 215102 492938 234546 493174
rect 234782 492938 234866 493174
rect 235102 492938 254546 493174
rect 254782 492938 254866 493174
rect 255102 492938 274546 493174
rect 274782 492938 274866 493174
rect 275102 492938 294546 493174
rect 294782 492938 294866 493174
rect 295102 492938 314546 493174
rect 314782 492938 314866 493174
rect 315102 492938 334546 493174
rect 334782 492938 334866 493174
rect 335102 492938 354546 493174
rect 354782 492938 354866 493174
rect 355102 492938 374546 493174
rect 374782 492938 374866 493174
rect 375102 492938 394546 493174
rect 394782 492938 394866 493174
rect 395102 492938 414546 493174
rect 414782 492938 414866 493174
rect 415102 492938 434546 493174
rect 434782 492938 434866 493174
rect 435102 492938 454546 493174
rect 454782 492938 454866 493174
rect 455102 492938 474546 493174
rect 474782 492938 474866 493174
rect 475102 492938 494546 493174
rect 494782 492938 494866 493174
rect 495102 492938 514546 493174
rect 514782 492938 514866 493174
rect 515102 492938 534546 493174
rect 534782 492938 534866 493174
rect 535102 492938 554546 493174
rect 554782 492938 554866 493174
rect 555102 492938 574546 493174
rect 574782 492938 574866 493174
rect 575102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 14546 492854
rect 14782 492618 14866 492854
rect 15102 492618 34546 492854
rect 34782 492618 34866 492854
rect 35102 492618 54546 492854
rect 54782 492618 54866 492854
rect 55102 492618 74546 492854
rect 74782 492618 74866 492854
rect 75102 492618 94546 492854
rect 94782 492618 94866 492854
rect 95102 492618 114546 492854
rect 114782 492618 114866 492854
rect 115102 492618 134546 492854
rect 134782 492618 134866 492854
rect 135102 492618 154546 492854
rect 154782 492618 154866 492854
rect 155102 492618 174546 492854
rect 174782 492618 174866 492854
rect 175102 492618 194546 492854
rect 194782 492618 194866 492854
rect 195102 492618 214546 492854
rect 214782 492618 214866 492854
rect 215102 492618 234546 492854
rect 234782 492618 234866 492854
rect 235102 492618 254546 492854
rect 254782 492618 254866 492854
rect 255102 492618 274546 492854
rect 274782 492618 274866 492854
rect 275102 492618 294546 492854
rect 294782 492618 294866 492854
rect 295102 492618 314546 492854
rect 314782 492618 314866 492854
rect 315102 492618 334546 492854
rect 334782 492618 334866 492854
rect 335102 492618 354546 492854
rect 354782 492618 354866 492854
rect 355102 492618 374546 492854
rect 374782 492618 374866 492854
rect 375102 492618 394546 492854
rect 394782 492618 394866 492854
rect 395102 492618 414546 492854
rect 414782 492618 414866 492854
rect 415102 492618 434546 492854
rect 434782 492618 434866 492854
rect 435102 492618 454546 492854
rect 454782 492618 454866 492854
rect 455102 492618 474546 492854
rect 474782 492618 474866 492854
rect 475102 492618 494546 492854
rect 494782 492618 494866 492854
rect 495102 492618 514546 492854
rect 514782 492618 514866 492854
rect 515102 492618 534546 492854
rect 534782 492618 534866 492854
rect 535102 492618 554546 492854
rect 554782 492618 554866 492854
rect 555102 492618 574546 492854
rect 574782 492618 574866 492854
rect 575102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 10826 489454
rect 11062 489218 11146 489454
rect 11382 489218 30826 489454
rect 31062 489218 31146 489454
rect 31382 489218 50826 489454
rect 51062 489218 51146 489454
rect 51382 489218 70826 489454
rect 71062 489218 71146 489454
rect 71382 489218 90826 489454
rect 91062 489218 91146 489454
rect 91382 489218 110826 489454
rect 111062 489218 111146 489454
rect 111382 489218 130826 489454
rect 131062 489218 131146 489454
rect 131382 489218 150826 489454
rect 151062 489218 151146 489454
rect 151382 489218 170826 489454
rect 171062 489218 171146 489454
rect 171382 489218 190826 489454
rect 191062 489218 191146 489454
rect 191382 489218 210826 489454
rect 211062 489218 211146 489454
rect 211382 489218 230826 489454
rect 231062 489218 231146 489454
rect 231382 489218 250826 489454
rect 251062 489218 251146 489454
rect 251382 489218 270826 489454
rect 271062 489218 271146 489454
rect 271382 489218 290826 489454
rect 291062 489218 291146 489454
rect 291382 489218 310826 489454
rect 311062 489218 311146 489454
rect 311382 489218 330826 489454
rect 331062 489218 331146 489454
rect 331382 489218 350826 489454
rect 351062 489218 351146 489454
rect 351382 489218 370826 489454
rect 371062 489218 371146 489454
rect 371382 489218 390826 489454
rect 391062 489218 391146 489454
rect 391382 489218 410826 489454
rect 411062 489218 411146 489454
rect 411382 489218 430826 489454
rect 431062 489218 431146 489454
rect 431382 489218 450826 489454
rect 451062 489218 451146 489454
rect 451382 489218 470826 489454
rect 471062 489218 471146 489454
rect 471382 489218 490826 489454
rect 491062 489218 491146 489454
rect 491382 489218 510826 489454
rect 511062 489218 511146 489454
rect 511382 489218 530826 489454
rect 531062 489218 531146 489454
rect 531382 489218 550826 489454
rect 551062 489218 551146 489454
rect 551382 489218 570826 489454
rect 571062 489218 571146 489454
rect 571382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 10826 489134
rect 11062 488898 11146 489134
rect 11382 488898 30826 489134
rect 31062 488898 31146 489134
rect 31382 488898 50826 489134
rect 51062 488898 51146 489134
rect 51382 488898 70826 489134
rect 71062 488898 71146 489134
rect 71382 488898 90826 489134
rect 91062 488898 91146 489134
rect 91382 488898 110826 489134
rect 111062 488898 111146 489134
rect 111382 488898 130826 489134
rect 131062 488898 131146 489134
rect 131382 488898 150826 489134
rect 151062 488898 151146 489134
rect 151382 488898 170826 489134
rect 171062 488898 171146 489134
rect 171382 488898 190826 489134
rect 191062 488898 191146 489134
rect 191382 488898 210826 489134
rect 211062 488898 211146 489134
rect 211382 488898 230826 489134
rect 231062 488898 231146 489134
rect 231382 488898 250826 489134
rect 251062 488898 251146 489134
rect 251382 488898 270826 489134
rect 271062 488898 271146 489134
rect 271382 488898 290826 489134
rect 291062 488898 291146 489134
rect 291382 488898 310826 489134
rect 311062 488898 311146 489134
rect 311382 488898 330826 489134
rect 331062 488898 331146 489134
rect 331382 488898 350826 489134
rect 351062 488898 351146 489134
rect 351382 488898 370826 489134
rect 371062 488898 371146 489134
rect 371382 488898 390826 489134
rect 391062 488898 391146 489134
rect 391382 488898 410826 489134
rect 411062 488898 411146 489134
rect 411382 488898 430826 489134
rect 431062 488898 431146 489134
rect 431382 488898 450826 489134
rect 451062 488898 451146 489134
rect 451382 488898 470826 489134
rect 471062 488898 471146 489134
rect 471382 488898 490826 489134
rect 491062 488898 491146 489134
rect 491382 488898 510826 489134
rect 511062 488898 511146 489134
rect 511382 488898 530826 489134
rect 531062 488898 531146 489134
rect 531382 488898 550826 489134
rect 551062 488898 551146 489134
rect 551382 488898 570826 489134
rect 571062 488898 571146 489134
rect 571382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 11986 482614
rect 12222 482378 12306 482614
rect 12542 482378 31986 482614
rect 32222 482378 32306 482614
rect 32542 482378 51986 482614
rect 52222 482378 52306 482614
rect 52542 482378 71986 482614
rect 72222 482378 72306 482614
rect 72542 482378 91986 482614
rect 92222 482378 92306 482614
rect 92542 482378 111986 482614
rect 112222 482378 112306 482614
rect 112542 482378 131986 482614
rect 132222 482378 132306 482614
rect 132542 482378 151986 482614
rect 152222 482378 152306 482614
rect 152542 482378 171986 482614
rect 172222 482378 172306 482614
rect 172542 482378 191986 482614
rect 192222 482378 192306 482614
rect 192542 482378 211986 482614
rect 212222 482378 212306 482614
rect 212542 482378 231986 482614
rect 232222 482378 232306 482614
rect 232542 482378 251986 482614
rect 252222 482378 252306 482614
rect 252542 482378 271986 482614
rect 272222 482378 272306 482614
rect 272542 482378 291986 482614
rect 292222 482378 292306 482614
rect 292542 482378 311986 482614
rect 312222 482378 312306 482614
rect 312542 482378 331986 482614
rect 332222 482378 332306 482614
rect 332542 482378 351986 482614
rect 352222 482378 352306 482614
rect 352542 482378 371986 482614
rect 372222 482378 372306 482614
rect 372542 482378 391986 482614
rect 392222 482378 392306 482614
rect 392542 482378 411986 482614
rect 412222 482378 412306 482614
rect 412542 482378 431986 482614
rect 432222 482378 432306 482614
rect 432542 482378 451986 482614
rect 452222 482378 452306 482614
rect 452542 482378 471986 482614
rect 472222 482378 472306 482614
rect 472542 482378 491986 482614
rect 492222 482378 492306 482614
rect 492542 482378 511986 482614
rect 512222 482378 512306 482614
rect 512542 482378 531986 482614
rect 532222 482378 532306 482614
rect 532542 482378 551986 482614
rect 552222 482378 552306 482614
rect 552542 482378 571986 482614
rect 572222 482378 572306 482614
rect 572542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 11986 482294
rect 12222 482058 12306 482294
rect 12542 482058 31986 482294
rect 32222 482058 32306 482294
rect 32542 482058 51986 482294
rect 52222 482058 52306 482294
rect 52542 482058 71986 482294
rect 72222 482058 72306 482294
rect 72542 482058 91986 482294
rect 92222 482058 92306 482294
rect 92542 482058 111986 482294
rect 112222 482058 112306 482294
rect 112542 482058 131986 482294
rect 132222 482058 132306 482294
rect 132542 482058 151986 482294
rect 152222 482058 152306 482294
rect 152542 482058 171986 482294
rect 172222 482058 172306 482294
rect 172542 482058 191986 482294
rect 192222 482058 192306 482294
rect 192542 482058 211986 482294
rect 212222 482058 212306 482294
rect 212542 482058 231986 482294
rect 232222 482058 232306 482294
rect 232542 482058 251986 482294
rect 252222 482058 252306 482294
rect 252542 482058 271986 482294
rect 272222 482058 272306 482294
rect 272542 482058 291986 482294
rect 292222 482058 292306 482294
rect 292542 482058 311986 482294
rect 312222 482058 312306 482294
rect 312542 482058 331986 482294
rect 332222 482058 332306 482294
rect 332542 482058 351986 482294
rect 352222 482058 352306 482294
rect 352542 482058 371986 482294
rect 372222 482058 372306 482294
rect 372542 482058 391986 482294
rect 392222 482058 392306 482294
rect 392542 482058 411986 482294
rect 412222 482058 412306 482294
rect 412542 482058 431986 482294
rect 432222 482058 432306 482294
rect 432542 482058 451986 482294
rect 452222 482058 452306 482294
rect 452542 482058 471986 482294
rect 472222 482058 472306 482294
rect 472542 482058 491986 482294
rect 492222 482058 492306 482294
rect 492542 482058 511986 482294
rect 512222 482058 512306 482294
rect 512542 482058 531986 482294
rect 532222 482058 532306 482294
rect 532542 482058 551986 482294
rect 552222 482058 552306 482294
rect 552542 482058 571986 482294
rect 572222 482058 572306 482294
rect 572542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 8266 478894
rect 8502 478658 8586 478894
rect 8822 478658 28266 478894
rect 28502 478658 28586 478894
rect 28822 478658 48266 478894
rect 48502 478658 48586 478894
rect 48822 478658 68266 478894
rect 68502 478658 68586 478894
rect 68822 478658 88266 478894
rect 88502 478658 88586 478894
rect 88822 478658 108266 478894
rect 108502 478658 108586 478894
rect 108822 478658 128266 478894
rect 128502 478658 128586 478894
rect 128822 478658 148266 478894
rect 148502 478658 148586 478894
rect 148822 478658 168266 478894
rect 168502 478658 168586 478894
rect 168822 478658 188266 478894
rect 188502 478658 188586 478894
rect 188822 478658 208266 478894
rect 208502 478658 208586 478894
rect 208822 478658 228266 478894
rect 228502 478658 228586 478894
rect 228822 478658 248266 478894
rect 248502 478658 248586 478894
rect 248822 478658 268266 478894
rect 268502 478658 268586 478894
rect 268822 478658 288266 478894
rect 288502 478658 288586 478894
rect 288822 478658 308266 478894
rect 308502 478658 308586 478894
rect 308822 478658 328266 478894
rect 328502 478658 328586 478894
rect 328822 478658 348266 478894
rect 348502 478658 348586 478894
rect 348822 478658 368266 478894
rect 368502 478658 368586 478894
rect 368822 478658 388266 478894
rect 388502 478658 388586 478894
rect 388822 478658 408266 478894
rect 408502 478658 408586 478894
rect 408822 478658 428266 478894
rect 428502 478658 428586 478894
rect 428822 478658 448266 478894
rect 448502 478658 448586 478894
rect 448822 478658 468266 478894
rect 468502 478658 468586 478894
rect 468822 478658 488266 478894
rect 488502 478658 488586 478894
rect 488822 478658 508266 478894
rect 508502 478658 508586 478894
rect 508822 478658 528266 478894
rect 528502 478658 528586 478894
rect 528822 478658 548266 478894
rect 548502 478658 548586 478894
rect 548822 478658 568266 478894
rect 568502 478658 568586 478894
rect 568822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 8266 478574
rect 8502 478338 8586 478574
rect 8822 478338 28266 478574
rect 28502 478338 28586 478574
rect 28822 478338 48266 478574
rect 48502 478338 48586 478574
rect 48822 478338 68266 478574
rect 68502 478338 68586 478574
rect 68822 478338 88266 478574
rect 88502 478338 88586 478574
rect 88822 478338 108266 478574
rect 108502 478338 108586 478574
rect 108822 478338 128266 478574
rect 128502 478338 128586 478574
rect 128822 478338 148266 478574
rect 148502 478338 148586 478574
rect 148822 478338 168266 478574
rect 168502 478338 168586 478574
rect 168822 478338 188266 478574
rect 188502 478338 188586 478574
rect 188822 478338 208266 478574
rect 208502 478338 208586 478574
rect 208822 478338 228266 478574
rect 228502 478338 228586 478574
rect 228822 478338 248266 478574
rect 248502 478338 248586 478574
rect 248822 478338 268266 478574
rect 268502 478338 268586 478574
rect 268822 478338 288266 478574
rect 288502 478338 288586 478574
rect 288822 478338 308266 478574
rect 308502 478338 308586 478574
rect 308822 478338 328266 478574
rect 328502 478338 328586 478574
rect 328822 478338 348266 478574
rect 348502 478338 348586 478574
rect 348822 478338 368266 478574
rect 368502 478338 368586 478574
rect 368822 478338 388266 478574
rect 388502 478338 388586 478574
rect 388822 478338 408266 478574
rect 408502 478338 408586 478574
rect 408822 478338 428266 478574
rect 428502 478338 428586 478574
rect 428822 478338 448266 478574
rect 448502 478338 448586 478574
rect 448822 478338 468266 478574
rect 468502 478338 468586 478574
rect 468822 478338 488266 478574
rect 488502 478338 488586 478574
rect 488822 478338 508266 478574
rect 508502 478338 508586 478574
rect 508822 478338 528266 478574
rect 528502 478338 528586 478574
rect 528822 478338 548266 478574
rect 548502 478338 548586 478574
rect 548822 478338 568266 478574
rect 568502 478338 568586 478574
rect 568822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 4546 475174
rect 4782 474938 4866 475174
rect 5102 474938 24546 475174
rect 24782 474938 24866 475174
rect 25102 474938 44546 475174
rect 44782 474938 44866 475174
rect 45102 474938 64546 475174
rect 64782 474938 64866 475174
rect 65102 474938 84546 475174
rect 84782 474938 84866 475174
rect 85102 474938 104546 475174
rect 104782 474938 104866 475174
rect 105102 474938 124546 475174
rect 124782 474938 124866 475174
rect 125102 474938 144546 475174
rect 144782 474938 144866 475174
rect 145102 474938 164546 475174
rect 164782 474938 164866 475174
rect 165102 474938 184546 475174
rect 184782 474938 184866 475174
rect 185102 474938 204546 475174
rect 204782 474938 204866 475174
rect 205102 474938 224546 475174
rect 224782 474938 224866 475174
rect 225102 474938 244546 475174
rect 244782 474938 244866 475174
rect 245102 474938 264546 475174
rect 264782 474938 264866 475174
rect 265102 474938 284546 475174
rect 284782 474938 284866 475174
rect 285102 474938 304546 475174
rect 304782 474938 304866 475174
rect 305102 474938 324546 475174
rect 324782 474938 324866 475174
rect 325102 474938 344546 475174
rect 344782 474938 344866 475174
rect 345102 474938 364546 475174
rect 364782 474938 364866 475174
rect 365102 474938 384546 475174
rect 384782 474938 384866 475174
rect 385102 474938 404546 475174
rect 404782 474938 404866 475174
rect 405102 474938 424546 475174
rect 424782 474938 424866 475174
rect 425102 474938 444546 475174
rect 444782 474938 444866 475174
rect 445102 474938 464546 475174
rect 464782 474938 464866 475174
rect 465102 474938 484546 475174
rect 484782 474938 484866 475174
rect 485102 474938 504546 475174
rect 504782 474938 504866 475174
rect 505102 474938 524546 475174
rect 524782 474938 524866 475174
rect 525102 474938 544546 475174
rect 544782 474938 544866 475174
rect 545102 474938 564546 475174
rect 564782 474938 564866 475174
rect 565102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 4546 474854
rect 4782 474618 4866 474854
rect 5102 474618 24546 474854
rect 24782 474618 24866 474854
rect 25102 474618 44546 474854
rect 44782 474618 44866 474854
rect 45102 474618 64546 474854
rect 64782 474618 64866 474854
rect 65102 474618 84546 474854
rect 84782 474618 84866 474854
rect 85102 474618 104546 474854
rect 104782 474618 104866 474854
rect 105102 474618 124546 474854
rect 124782 474618 124866 474854
rect 125102 474618 144546 474854
rect 144782 474618 144866 474854
rect 145102 474618 164546 474854
rect 164782 474618 164866 474854
rect 165102 474618 184546 474854
rect 184782 474618 184866 474854
rect 185102 474618 204546 474854
rect 204782 474618 204866 474854
rect 205102 474618 224546 474854
rect 224782 474618 224866 474854
rect 225102 474618 244546 474854
rect 244782 474618 244866 474854
rect 245102 474618 264546 474854
rect 264782 474618 264866 474854
rect 265102 474618 284546 474854
rect 284782 474618 284866 474854
rect 285102 474618 304546 474854
rect 304782 474618 304866 474854
rect 305102 474618 324546 474854
rect 324782 474618 324866 474854
rect 325102 474618 344546 474854
rect 344782 474618 344866 474854
rect 345102 474618 364546 474854
rect 364782 474618 364866 474854
rect 365102 474618 384546 474854
rect 384782 474618 384866 474854
rect 385102 474618 404546 474854
rect 404782 474618 404866 474854
rect 405102 474618 424546 474854
rect 424782 474618 424866 474854
rect 425102 474618 444546 474854
rect 444782 474618 444866 474854
rect 445102 474618 464546 474854
rect 464782 474618 464866 474854
rect 465102 474618 484546 474854
rect 484782 474618 484866 474854
rect 485102 474618 504546 474854
rect 504782 474618 504866 474854
rect 505102 474618 524546 474854
rect 524782 474618 524866 474854
rect 525102 474618 544546 474854
rect 544782 474618 544866 474854
rect 545102 474618 564546 474854
rect 564782 474618 564866 474854
rect 565102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 826 471454
rect 1062 471218 1146 471454
rect 1382 471218 20826 471454
rect 21062 471218 21146 471454
rect 21382 471218 40826 471454
rect 41062 471218 41146 471454
rect 41382 471218 60826 471454
rect 61062 471218 61146 471454
rect 61382 471218 80826 471454
rect 81062 471218 81146 471454
rect 81382 471218 100826 471454
rect 101062 471218 101146 471454
rect 101382 471218 120826 471454
rect 121062 471218 121146 471454
rect 121382 471218 140826 471454
rect 141062 471218 141146 471454
rect 141382 471218 160826 471454
rect 161062 471218 161146 471454
rect 161382 471218 180826 471454
rect 181062 471218 181146 471454
rect 181382 471218 200826 471454
rect 201062 471218 201146 471454
rect 201382 471218 220826 471454
rect 221062 471218 221146 471454
rect 221382 471218 240826 471454
rect 241062 471218 241146 471454
rect 241382 471218 260826 471454
rect 261062 471218 261146 471454
rect 261382 471218 280826 471454
rect 281062 471218 281146 471454
rect 281382 471218 300826 471454
rect 301062 471218 301146 471454
rect 301382 471218 320826 471454
rect 321062 471218 321146 471454
rect 321382 471218 340826 471454
rect 341062 471218 341146 471454
rect 341382 471218 360826 471454
rect 361062 471218 361146 471454
rect 361382 471218 380826 471454
rect 381062 471218 381146 471454
rect 381382 471218 400826 471454
rect 401062 471218 401146 471454
rect 401382 471218 420826 471454
rect 421062 471218 421146 471454
rect 421382 471218 440826 471454
rect 441062 471218 441146 471454
rect 441382 471218 460826 471454
rect 461062 471218 461146 471454
rect 461382 471218 480826 471454
rect 481062 471218 481146 471454
rect 481382 471218 500826 471454
rect 501062 471218 501146 471454
rect 501382 471218 520826 471454
rect 521062 471218 521146 471454
rect 521382 471218 540826 471454
rect 541062 471218 541146 471454
rect 541382 471218 560826 471454
rect 561062 471218 561146 471454
rect 561382 471218 580826 471454
rect 581062 471218 581146 471454
rect 581382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 826 471134
rect 1062 470898 1146 471134
rect 1382 470898 20826 471134
rect 21062 470898 21146 471134
rect 21382 470898 40826 471134
rect 41062 470898 41146 471134
rect 41382 470898 60826 471134
rect 61062 470898 61146 471134
rect 61382 470898 80826 471134
rect 81062 470898 81146 471134
rect 81382 470898 100826 471134
rect 101062 470898 101146 471134
rect 101382 470898 120826 471134
rect 121062 470898 121146 471134
rect 121382 470898 140826 471134
rect 141062 470898 141146 471134
rect 141382 470898 160826 471134
rect 161062 470898 161146 471134
rect 161382 470898 180826 471134
rect 181062 470898 181146 471134
rect 181382 470898 200826 471134
rect 201062 470898 201146 471134
rect 201382 470898 220826 471134
rect 221062 470898 221146 471134
rect 221382 470898 240826 471134
rect 241062 470898 241146 471134
rect 241382 470898 260826 471134
rect 261062 470898 261146 471134
rect 261382 470898 280826 471134
rect 281062 470898 281146 471134
rect 281382 470898 300826 471134
rect 301062 470898 301146 471134
rect 301382 470898 320826 471134
rect 321062 470898 321146 471134
rect 321382 470898 340826 471134
rect 341062 470898 341146 471134
rect 341382 470898 360826 471134
rect 361062 470898 361146 471134
rect 361382 470898 380826 471134
rect 381062 470898 381146 471134
rect 381382 470898 400826 471134
rect 401062 470898 401146 471134
rect 401382 470898 420826 471134
rect 421062 470898 421146 471134
rect 421382 470898 440826 471134
rect 441062 470898 441146 471134
rect 441382 470898 460826 471134
rect 461062 470898 461146 471134
rect 461382 470898 480826 471134
rect 481062 470898 481146 471134
rect 481382 470898 500826 471134
rect 501062 470898 501146 471134
rect 501382 470898 520826 471134
rect 521062 470898 521146 471134
rect 521382 470898 540826 471134
rect 541062 470898 541146 471134
rect 541382 470898 560826 471134
rect 561062 470898 561146 471134
rect 561382 470898 580826 471134
rect 581062 470898 581146 471134
rect 581382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 21986 464614
rect 22222 464378 22306 464614
rect 22542 464378 41986 464614
rect 42222 464378 42306 464614
rect 42542 464378 61986 464614
rect 62222 464378 62306 464614
rect 62542 464378 81986 464614
rect 82222 464378 82306 464614
rect 82542 464378 101986 464614
rect 102222 464378 102306 464614
rect 102542 464378 121986 464614
rect 122222 464378 122306 464614
rect 122542 464378 141986 464614
rect 142222 464378 142306 464614
rect 142542 464378 161986 464614
rect 162222 464378 162306 464614
rect 162542 464378 181986 464614
rect 182222 464378 182306 464614
rect 182542 464378 201986 464614
rect 202222 464378 202306 464614
rect 202542 464378 221986 464614
rect 222222 464378 222306 464614
rect 222542 464378 241986 464614
rect 242222 464378 242306 464614
rect 242542 464378 261986 464614
rect 262222 464378 262306 464614
rect 262542 464378 281986 464614
rect 282222 464378 282306 464614
rect 282542 464378 301986 464614
rect 302222 464378 302306 464614
rect 302542 464378 321986 464614
rect 322222 464378 322306 464614
rect 322542 464378 341986 464614
rect 342222 464378 342306 464614
rect 342542 464378 361986 464614
rect 362222 464378 362306 464614
rect 362542 464378 381986 464614
rect 382222 464378 382306 464614
rect 382542 464378 401986 464614
rect 402222 464378 402306 464614
rect 402542 464378 421986 464614
rect 422222 464378 422306 464614
rect 422542 464378 441986 464614
rect 442222 464378 442306 464614
rect 442542 464378 461986 464614
rect 462222 464378 462306 464614
rect 462542 464378 481986 464614
rect 482222 464378 482306 464614
rect 482542 464378 501986 464614
rect 502222 464378 502306 464614
rect 502542 464378 521986 464614
rect 522222 464378 522306 464614
rect 522542 464378 541986 464614
rect 542222 464378 542306 464614
rect 542542 464378 561986 464614
rect 562222 464378 562306 464614
rect 562542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 21986 464294
rect 22222 464058 22306 464294
rect 22542 464058 41986 464294
rect 42222 464058 42306 464294
rect 42542 464058 61986 464294
rect 62222 464058 62306 464294
rect 62542 464058 81986 464294
rect 82222 464058 82306 464294
rect 82542 464058 101986 464294
rect 102222 464058 102306 464294
rect 102542 464058 121986 464294
rect 122222 464058 122306 464294
rect 122542 464058 141986 464294
rect 142222 464058 142306 464294
rect 142542 464058 161986 464294
rect 162222 464058 162306 464294
rect 162542 464058 181986 464294
rect 182222 464058 182306 464294
rect 182542 464058 201986 464294
rect 202222 464058 202306 464294
rect 202542 464058 221986 464294
rect 222222 464058 222306 464294
rect 222542 464058 241986 464294
rect 242222 464058 242306 464294
rect 242542 464058 261986 464294
rect 262222 464058 262306 464294
rect 262542 464058 281986 464294
rect 282222 464058 282306 464294
rect 282542 464058 301986 464294
rect 302222 464058 302306 464294
rect 302542 464058 321986 464294
rect 322222 464058 322306 464294
rect 322542 464058 341986 464294
rect 342222 464058 342306 464294
rect 342542 464058 361986 464294
rect 362222 464058 362306 464294
rect 362542 464058 381986 464294
rect 382222 464058 382306 464294
rect 382542 464058 401986 464294
rect 402222 464058 402306 464294
rect 402542 464058 421986 464294
rect 422222 464058 422306 464294
rect 422542 464058 441986 464294
rect 442222 464058 442306 464294
rect 442542 464058 461986 464294
rect 462222 464058 462306 464294
rect 462542 464058 481986 464294
rect 482222 464058 482306 464294
rect 482542 464058 501986 464294
rect 502222 464058 502306 464294
rect 502542 464058 521986 464294
rect 522222 464058 522306 464294
rect 522542 464058 541986 464294
rect 542222 464058 542306 464294
rect 542542 464058 561986 464294
rect 562222 464058 562306 464294
rect 562542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 18266 460894
rect 18502 460658 18586 460894
rect 18822 460658 38266 460894
rect 38502 460658 38586 460894
rect 38822 460658 58266 460894
rect 58502 460658 58586 460894
rect 58822 460658 78266 460894
rect 78502 460658 78586 460894
rect 78822 460658 98266 460894
rect 98502 460658 98586 460894
rect 98822 460658 118266 460894
rect 118502 460658 118586 460894
rect 118822 460658 138266 460894
rect 138502 460658 138586 460894
rect 138822 460658 158266 460894
rect 158502 460658 158586 460894
rect 158822 460658 178266 460894
rect 178502 460658 178586 460894
rect 178822 460658 198266 460894
rect 198502 460658 198586 460894
rect 198822 460658 218266 460894
rect 218502 460658 218586 460894
rect 218822 460658 238266 460894
rect 238502 460658 238586 460894
rect 238822 460658 258266 460894
rect 258502 460658 258586 460894
rect 258822 460658 278266 460894
rect 278502 460658 278586 460894
rect 278822 460658 298266 460894
rect 298502 460658 298586 460894
rect 298822 460658 318266 460894
rect 318502 460658 318586 460894
rect 318822 460658 338266 460894
rect 338502 460658 338586 460894
rect 338822 460658 358266 460894
rect 358502 460658 358586 460894
rect 358822 460658 378266 460894
rect 378502 460658 378586 460894
rect 378822 460658 398266 460894
rect 398502 460658 398586 460894
rect 398822 460658 418266 460894
rect 418502 460658 418586 460894
rect 418822 460658 438266 460894
rect 438502 460658 438586 460894
rect 438822 460658 458266 460894
rect 458502 460658 458586 460894
rect 458822 460658 478266 460894
rect 478502 460658 478586 460894
rect 478822 460658 498266 460894
rect 498502 460658 498586 460894
rect 498822 460658 518266 460894
rect 518502 460658 518586 460894
rect 518822 460658 538266 460894
rect 538502 460658 538586 460894
rect 538822 460658 558266 460894
rect 558502 460658 558586 460894
rect 558822 460658 578266 460894
rect 578502 460658 578586 460894
rect 578822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 18266 460574
rect 18502 460338 18586 460574
rect 18822 460338 38266 460574
rect 38502 460338 38586 460574
rect 38822 460338 58266 460574
rect 58502 460338 58586 460574
rect 58822 460338 78266 460574
rect 78502 460338 78586 460574
rect 78822 460338 98266 460574
rect 98502 460338 98586 460574
rect 98822 460338 118266 460574
rect 118502 460338 118586 460574
rect 118822 460338 138266 460574
rect 138502 460338 138586 460574
rect 138822 460338 158266 460574
rect 158502 460338 158586 460574
rect 158822 460338 178266 460574
rect 178502 460338 178586 460574
rect 178822 460338 198266 460574
rect 198502 460338 198586 460574
rect 198822 460338 218266 460574
rect 218502 460338 218586 460574
rect 218822 460338 238266 460574
rect 238502 460338 238586 460574
rect 238822 460338 258266 460574
rect 258502 460338 258586 460574
rect 258822 460338 278266 460574
rect 278502 460338 278586 460574
rect 278822 460338 298266 460574
rect 298502 460338 298586 460574
rect 298822 460338 318266 460574
rect 318502 460338 318586 460574
rect 318822 460338 338266 460574
rect 338502 460338 338586 460574
rect 338822 460338 358266 460574
rect 358502 460338 358586 460574
rect 358822 460338 378266 460574
rect 378502 460338 378586 460574
rect 378822 460338 398266 460574
rect 398502 460338 398586 460574
rect 398822 460338 418266 460574
rect 418502 460338 418586 460574
rect 418822 460338 438266 460574
rect 438502 460338 438586 460574
rect 438822 460338 458266 460574
rect 458502 460338 458586 460574
rect 458822 460338 478266 460574
rect 478502 460338 478586 460574
rect 478822 460338 498266 460574
rect 498502 460338 498586 460574
rect 498822 460338 518266 460574
rect 518502 460338 518586 460574
rect 518822 460338 538266 460574
rect 538502 460338 538586 460574
rect 538822 460338 558266 460574
rect 558502 460338 558586 460574
rect 558822 460338 578266 460574
rect 578502 460338 578586 460574
rect 578822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 14546 457174
rect 14782 456938 14866 457174
rect 15102 456938 34546 457174
rect 34782 456938 34866 457174
rect 35102 456938 54546 457174
rect 54782 456938 54866 457174
rect 55102 456938 74546 457174
rect 74782 456938 74866 457174
rect 75102 456938 94546 457174
rect 94782 456938 94866 457174
rect 95102 456938 114546 457174
rect 114782 456938 114866 457174
rect 115102 456938 134546 457174
rect 134782 456938 134866 457174
rect 135102 456938 154546 457174
rect 154782 456938 154866 457174
rect 155102 456938 174546 457174
rect 174782 456938 174866 457174
rect 175102 456938 194546 457174
rect 194782 456938 194866 457174
rect 195102 456938 214546 457174
rect 214782 456938 214866 457174
rect 215102 456938 234546 457174
rect 234782 456938 234866 457174
rect 235102 456938 254546 457174
rect 254782 456938 254866 457174
rect 255102 456938 274546 457174
rect 274782 456938 274866 457174
rect 275102 456938 294546 457174
rect 294782 456938 294866 457174
rect 295102 456938 314546 457174
rect 314782 456938 314866 457174
rect 315102 456938 334546 457174
rect 334782 456938 334866 457174
rect 335102 456938 354546 457174
rect 354782 456938 354866 457174
rect 355102 456938 374546 457174
rect 374782 456938 374866 457174
rect 375102 456938 394546 457174
rect 394782 456938 394866 457174
rect 395102 456938 414546 457174
rect 414782 456938 414866 457174
rect 415102 456938 434546 457174
rect 434782 456938 434866 457174
rect 435102 456938 454546 457174
rect 454782 456938 454866 457174
rect 455102 456938 474546 457174
rect 474782 456938 474866 457174
rect 475102 456938 494546 457174
rect 494782 456938 494866 457174
rect 495102 456938 514546 457174
rect 514782 456938 514866 457174
rect 515102 456938 534546 457174
rect 534782 456938 534866 457174
rect 535102 456938 554546 457174
rect 554782 456938 554866 457174
rect 555102 456938 574546 457174
rect 574782 456938 574866 457174
rect 575102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 14546 456854
rect 14782 456618 14866 456854
rect 15102 456618 34546 456854
rect 34782 456618 34866 456854
rect 35102 456618 54546 456854
rect 54782 456618 54866 456854
rect 55102 456618 74546 456854
rect 74782 456618 74866 456854
rect 75102 456618 94546 456854
rect 94782 456618 94866 456854
rect 95102 456618 114546 456854
rect 114782 456618 114866 456854
rect 115102 456618 134546 456854
rect 134782 456618 134866 456854
rect 135102 456618 154546 456854
rect 154782 456618 154866 456854
rect 155102 456618 174546 456854
rect 174782 456618 174866 456854
rect 175102 456618 194546 456854
rect 194782 456618 194866 456854
rect 195102 456618 214546 456854
rect 214782 456618 214866 456854
rect 215102 456618 234546 456854
rect 234782 456618 234866 456854
rect 235102 456618 254546 456854
rect 254782 456618 254866 456854
rect 255102 456618 274546 456854
rect 274782 456618 274866 456854
rect 275102 456618 294546 456854
rect 294782 456618 294866 456854
rect 295102 456618 314546 456854
rect 314782 456618 314866 456854
rect 315102 456618 334546 456854
rect 334782 456618 334866 456854
rect 335102 456618 354546 456854
rect 354782 456618 354866 456854
rect 355102 456618 374546 456854
rect 374782 456618 374866 456854
rect 375102 456618 394546 456854
rect 394782 456618 394866 456854
rect 395102 456618 414546 456854
rect 414782 456618 414866 456854
rect 415102 456618 434546 456854
rect 434782 456618 434866 456854
rect 435102 456618 454546 456854
rect 454782 456618 454866 456854
rect 455102 456618 474546 456854
rect 474782 456618 474866 456854
rect 475102 456618 494546 456854
rect 494782 456618 494866 456854
rect 495102 456618 514546 456854
rect 514782 456618 514866 456854
rect 515102 456618 534546 456854
rect 534782 456618 534866 456854
rect 535102 456618 554546 456854
rect 554782 456618 554866 456854
rect 555102 456618 574546 456854
rect 574782 456618 574866 456854
rect 575102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 10826 453454
rect 11062 453218 11146 453454
rect 11382 453218 30826 453454
rect 31062 453218 31146 453454
rect 31382 453218 50826 453454
rect 51062 453218 51146 453454
rect 51382 453218 70826 453454
rect 71062 453218 71146 453454
rect 71382 453218 90826 453454
rect 91062 453218 91146 453454
rect 91382 453218 110826 453454
rect 111062 453218 111146 453454
rect 111382 453218 130826 453454
rect 131062 453218 131146 453454
rect 131382 453218 150826 453454
rect 151062 453218 151146 453454
rect 151382 453218 170826 453454
rect 171062 453218 171146 453454
rect 171382 453218 190826 453454
rect 191062 453218 191146 453454
rect 191382 453218 210826 453454
rect 211062 453218 211146 453454
rect 211382 453218 230826 453454
rect 231062 453218 231146 453454
rect 231382 453218 250826 453454
rect 251062 453218 251146 453454
rect 251382 453218 270826 453454
rect 271062 453218 271146 453454
rect 271382 453218 290826 453454
rect 291062 453218 291146 453454
rect 291382 453218 310826 453454
rect 311062 453218 311146 453454
rect 311382 453218 330826 453454
rect 331062 453218 331146 453454
rect 331382 453218 350826 453454
rect 351062 453218 351146 453454
rect 351382 453218 370826 453454
rect 371062 453218 371146 453454
rect 371382 453218 390826 453454
rect 391062 453218 391146 453454
rect 391382 453218 410826 453454
rect 411062 453218 411146 453454
rect 411382 453218 430826 453454
rect 431062 453218 431146 453454
rect 431382 453218 450826 453454
rect 451062 453218 451146 453454
rect 451382 453218 470826 453454
rect 471062 453218 471146 453454
rect 471382 453218 490826 453454
rect 491062 453218 491146 453454
rect 491382 453218 510826 453454
rect 511062 453218 511146 453454
rect 511382 453218 530826 453454
rect 531062 453218 531146 453454
rect 531382 453218 550826 453454
rect 551062 453218 551146 453454
rect 551382 453218 570826 453454
rect 571062 453218 571146 453454
rect 571382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 10826 453134
rect 11062 452898 11146 453134
rect 11382 452898 30826 453134
rect 31062 452898 31146 453134
rect 31382 452898 50826 453134
rect 51062 452898 51146 453134
rect 51382 452898 70826 453134
rect 71062 452898 71146 453134
rect 71382 452898 90826 453134
rect 91062 452898 91146 453134
rect 91382 452898 110826 453134
rect 111062 452898 111146 453134
rect 111382 452898 130826 453134
rect 131062 452898 131146 453134
rect 131382 452898 150826 453134
rect 151062 452898 151146 453134
rect 151382 452898 170826 453134
rect 171062 452898 171146 453134
rect 171382 452898 190826 453134
rect 191062 452898 191146 453134
rect 191382 452898 210826 453134
rect 211062 452898 211146 453134
rect 211382 452898 230826 453134
rect 231062 452898 231146 453134
rect 231382 452898 250826 453134
rect 251062 452898 251146 453134
rect 251382 452898 270826 453134
rect 271062 452898 271146 453134
rect 271382 452898 290826 453134
rect 291062 452898 291146 453134
rect 291382 452898 310826 453134
rect 311062 452898 311146 453134
rect 311382 452898 330826 453134
rect 331062 452898 331146 453134
rect 331382 452898 350826 453134
rect 351062 452898 351146 453134
rect 351382 452898 370826 453134
rect 371062 452898 371146 453134
rect 371382 452898 390826 453134
rect 391062 452898 391146 453134
rect 391382 452898 410826 453134
rect 411062 452898 411146 453134
rect 411382 452898 430826 453134
rect 431062 452898 431146 453134
rect 431382 452898 450826 453134
rect 451062 452898 451146 453134
rect 451382 452898 470826 453134
rect 471062 452898 471146 453134
rect 471382 452898 490826 453134
rect 491062 452898 491146 453134
rect 491382 452898 510826 453134
rect 511062 452898 511146 453134
rect 511382 452898 530826 453134
rect 531062 452898 531146 453134
rect 531382 452898 550826 453134
rect 551062 452898 551146 453134
rect 551382 452898 570826 453134
rect 571062 452898 571146 453134
rect 571382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 11986 446614
rect 12222 446378 12306 446614
rect 12542 446378 31986 446614
rect 32222 446378 32306 446614
rect 32542 446378 51986 446614
rect 52222 446378 52306 446614
rect 52542 446378 71986 446614
rect 72222 446378 72306 446614
rect 72542 446378 91986 446614
rect 92222 446378 92306 446614
rect 92542 446378 111986 446614
rect 112222 446378 112306 446614
rect 112542 446378 131986 446614
rect 132222 446378 132306 446614
rect 132542 446378 151986 446614
rect 152222 446378 152306 446614
rect 152542 446378 171986 446614
rect 172222 446378 172306 446614
rect 172542 446378 191986 446614
rect 192222 446378 192306 446614
rect 192542 446378 211986 446614
rect 212222 446378 212306 446614
rect 212542 446378 231986 446614
rect 232222 446378 232306 446614
rect 232542 446378 251986 446614
rect 252222 446378 252306 446614
rect 252542 446378 271986 446614
rect 272222 446378 272306 446614
rect 272542 446378 291986 446614
rect 292222 446378 292306 446614
rect 292542 446378 311986 446614
rect 312222 446378 312306 446614
rect 312542 446378 331986 446614
rect 332222 446378 332306 446614
rect 332542 446378 351986 446614
rect 352222 446378 352306 446614
rect 352542 446378 371986 446614
rect 372222 446378 372306 446614
rect 372542 446378 391986 446614
rect 392222 446378 392306 446614
rect 392542 446378 411986 446614
rect 412222 446378 412306 446614
rect 412542 446378 431986 446614
rect 432222 446378 432306 446614
rect 432542 446378 451986 446614
rect 452222 446378 452306 446614
rect 452542 446378 471986 446614
rect 472222 446378 472306 446614
rect 472542 446378 491986 446614
rect 492222 446378 492306 446614
rect 492542 446378 511986 446614
rect 512222 446378 512306 446614
rect 512542 446378 531986 446614
rect 532222 446378 532306 446614
rect 532542 446378 551986 446614
rect 552222 446378 552306 446614
rect 552542 446378 571986 446614
rect 572222 446378 572306 446614
rect 572542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 11986 446294
rect 12222 446058 12306 446294
rect 12542 446058 31986 446294
rect 32222 446058 32306 446294
rect 32542 446058 51986 446294
rect 52222 446058 52306 446294
rect 52542 446058 71986 446294
rect 72222 446058 72306 446294
rect 72542 446058 91986 446294
rect 92222 446058 92306 446294
rect 92542 446058 111986 446294
rect 112222 446058 112306 446294
rect 112542 446058 131986 446294
rect 132222 446058 132306 446294
rect 132542 446058 151986 446294
rect 152222 446058 152306 446294
rect 152542 446058 171986 446294
rect 172222 446058 172306 446294
rect 172542 446058 191986 446294
rect 192222 446058 192306 446294
rect 192542 446058 211986 446294
rect 212222 446058 212306 446294
rect 212542 446058 231986 446294
rect 232222 446058 232306 446294
rect 232542 446058 251986 446294
rect 252222 446058 252306 446294
rect 252542 446058 271986 446294
rect 272222 446058 272306 446294
rect 272542 446058 291986 446294
rect 292222 446058 292306 446294
rect 292542 446058 311986 446294
rect 312222 446058 312306 446294
rect 312542 446058 331986 446294
rect 332222 446058 332306 446294
rect 332542 446058 351986 446294
rect 352222 446058 352306 446294
rect 352542 446058 371986 446294
rect 372222 446058 372306 446294
rect 372542 446058 391986 446294
rect 392222 446058 392306 446294
rect 392542 446058 411986 446294
rect 412222 446058 412306 446294
rect 412542 446058 431986 446294
rect 432222 446058 432306 446294
rect 432542 446058 451986 446294
rect 452222 446058 452306 446294
rect 452542 446058 471986 446294
rect 472222 446058 472306 446294
rect 472542 446058 491986 446294
rect 492222 446058 492306 446294
rect 492542 446058 511986 446294
rect 512222 446058 512306 446294
rect 512542 446058 531986 446294
rect 532222 446058 532306 446294
rect 532542 446058 551986 446294
rect 552222 446058 552306 446294
rect 552542 446058 571986 446294
rect 572222 446058 572306 446294
rect 572542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 8266 442894
rect 8502 442658 8586 442894
rect 8822 442658 28266 442894
rect 28502 442658 28586 442894
rect 28822 442658 48266 442894
rect 48502 442658 48586 442894
rect 48822 442658 68266 442894
rect 68502 442658 68586 442894
rect 68822 442658 88266 442894
rect 88502 442658 88586 442894
rect 88822 442658 108266 442894
rect 108502 442658 108586 442894
rect 108822 442658 128266 442894
rect 128502 442658 128586 442894
rect 128822 442658 148266 442894
rect 148502 442658 148586 442894
rect 148822 442658 168266 442894
rect 168502 442658 168586 442894
rect 168822 442658 188266 442894
rect 188502 442658 188586 442894
rect 188822 442658 208266 442894
rect 208502 442658 208586 442894
rect 208822 442658 228266 442894
rect 228502 442658 228586 442894
rect 228822 442658 248266 442894
rect 248502 442658 248586 442894
rect 248822 442658 268266 442894
rect 268502 442658 268586 442894
rect 268822 442658 288266 442894
rect 288502 442658 288586 442894
rect 288822 442658 308266 442894
rect 308502 442658 308586 442894
rect 308822 442658 328266 442894
rect 328502 442658 328586 442894
rect 328822 442658 348266 442894
rect 348502 442658 348586 442894
rect 348822 442658 368266 442894
rect 368502 442658 368586 442894
rect 368822 442658 388266 442894
rect 388502 442658 388586 442894
rect 388822 442658 408266 442894
rect 408502 442658 408586 442894
rect 408822 442658 428266 442894
rect 428502 442658 428586 442894
rect 428822 442658 448266 442894
rect 448502 442658 448586 442894
rect 448822 442658 468266 442894
rect 468502 442658 468586 442894
rect 468822 442658 488266 442894
rect 488502 442658 488586 442894
rect 488822 442658 508266 442894
rect 508502 442658 508586 442894
rect 508822 442658 528266 442894
rect 528502 442658 528586 442894
rect 528822 442658 548266 442894
rect 548502 442658 548586 442894
rect 548822 442658 568266 442894
rect 568502 442658 568586 442894
rect 568822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 8266 442574
rect 8502 442338 8586 442574
rect 8822 442338 28266 442574
rect 28502 442338 28586 442574
rect 28822 442338 48266 442574
rect 48502 442338 48586 442574
rect 48822 442338 68266 442574
rect 68502 442338 68586 442574
rect 68822 442338 88266 442574
rect 88502 442338 88586 442574
rect 88822 442338 108266 442574
rect 108502 442338 108586 442574
rect 108822 442338 128266 442574
rect 128502 442338 128586 442574
rect 128822 442338 148266 442574
rect 148502 442338 148586 442574
rect 148822 442338 168266 442574
rect 168502 442338 168586 442574
rect 168822 442338 188266 442574
rect 188502 442338 188586 442574
rect 188822 442338 208266 442574
rect 208502 442338 208586 442574
rect 208822 442338 228266 442574
rect 228502 442338 228586 442574
rect 228822 442338 248266 442574
rect 248502 442338 248586 442574
rect 248822 442338 268266 442574
rect 268502 442338 268586 442574
rect 268822 442338 288266 442574
rect 288502 442338 288586 442574
rect 288822 442338 308266 442574
rect 308502 442338 308586 442574
rect 308822 442338 328266 442574
rect 328502 442338 328586 442574
rect 328822 442338 348266 442574
rect 348502 442338 348586 442574
rect 348822 442338 368266 442574
rect 368502 442338 368586 442574
rect 368822 442338 388266 442574
rect 388502 442338 388586 442574
rect 388822 442338 408266 442574
rect 408502 442338 408586 442574
rect 408822 442338 428266 442574
rect 428502 442338 428586 442574
rect 428822 442338 448266 442574
rect 448502 442338 448586 442574
rect 448822 442338 468266 442574
rect 468502 442338 468586 442574
rect 468822 442338 488266 442574
rect 488502 442338 488586 442574
rect 488822 442338 508266 442574
rect 508502 442338 508586 442574
rect 508822 442338 528266 442574
rect 528502 442338 528586 442574
rect 528822 442338 548266 442574
rect 548502 442338 548586 442574
rect 548822 442338 568266 442574
rect 568502 442338 568586 442574
rect 568822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 4546 439174
rect 4782 438938 4866 439174
rect 5102 438938 24546 439174
rect 24782 438938 24866 439174
rect 25102 438938 44546 439174
rect 44782 438938 44866 439174
rect 45102 438938 64546 439174
rect 64782 438938 64866 439174
rect 65102 438938 84546 439174
rect 84782 438938 84866 439174
rect 85102 438938 104546 439174
rect 104782 438938 104866 439174
rect 105102 438938 124546 439174
rect 124782 438938 124866 439174
rect 125102 438938 144546 439174
rect 144782 438938 144866 439174
rect 145102 438938 164546 439174
rect 164782 438938 164866 439174
rect 165102 438938 184546 439174
rect 184782 438938 184866 439174
rect 185102 438938 204546 439174
rect 204782 438938 204866 439174
rect 205102 438938 224546 439174
rect 224782 438938 224866 439174
rect 225102 438938 244546 439174
rect 244782 438938 244866 439174
rect 245102 438938 264546 439174
rect 264782 438938 264866 439174
rect 265102 438938 284546 439174
rect 284782 438938 284866 439174
rect 285102 438938 304546 439174
rect 304782 438938 304866 439174
rect 305102 438938 324546 439174
rect 324782 438938 324866 439174
rect 325102 438938 344546 439174
rect 344782 438938 344866 439174
rect 345102 438938 364546 439174
rect 364782 438938 364866 439174
rect 365102 438938 384546 439174
rect 384782 438938 384866 439174
rect 385102 438938 404546 439174
rect 404782 438938 404866 439174
rect 405102 438938 424546 439174
rect 424782 438938 424866 439174
rect 425102 438938 444546 439174
rect 444782 438938 444866 439174
rect 445102 438938 464546 439174
rect 464782 438938 464866 439174
rect 465102 438938 484546 439174
rect 484782 438938 484866 439174
rect 485102 438938 504546 439174
rect 504782 438938 504866 439174
rect 505102 438938 524546 439174
rect 524782 438938 524866 439174
rect 525102 438938 544546 439174
rect 544782 438938 544866 439174
rect 545102 438938 564546 439174
rect 564782 438938 564866 439174
rect 565102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 4546 438854
rect 4782 438618 4866 438854
rect 5102 438618 24546 438854
rect 24782 438618 24866 438854
rect 25102 438618 44546 438854
rect 44782 438618 44866 438854
rect 45102 438618 64546 438854
rect 64782 438618 64866 438854
rect 65102 438618 84546 438854
rect 84782 438618 84866 438854
rect 85102 438618 104546 438854
rect 104782 438618 104866 438854
rect 105102 438618 124546 438854
rect 124782 438618 124866 438854
rect 125102 438618 144546 438854
rect 144782 438618 144866 438854
rect 145102 438618 164546 438854
rect 164782 438618 164866 438854
rect 165102 438618 184546 438854
rect 184782 438618 184866 438854
rect 185102 438618 204546 438854
rect 204782 438618 204866 438854
rect 205102 438618 224546 438854
rect 224782 438618 224866 438854
rect 225102 438618 244546 438854
rect 244782 438618 244866 438854
rect 245102 438618 264546 438854
rect 264782 438618 264866 438854
rect 265102 438618 284546 438854
rect 284782 438618 284866 438854
rect 285102 438618 304546 438854
rect 304782 438618 304866 438854
rect 305102 438618 324546 438854
rect 324782 438618 324866 438854
rect 325102 438618 344546 438854
rect 344782 438618 344866 438854
rect 345102 438618 364546 438854
rect 364782 438618 364866 438854
rect 365102 438618 384546 438854
rect 384782 438618 384866 438854
rect 385102 438618 404546 438854
rect 404782 438618 404866 438854
rect 405102 438618 424546 438854
rect 424782 438618 424866 438854
rect 425102 438618 444546 438854
rect 444782 438618 444866 438854
rect 445102 438618 464546 438854
rect 464782 438618 464866 438854
rect 465102 438618 484546 438854
rect 484782 438618 484866 438854
rect 485102 438618 504546 438854
rect 504782 438618 504866 438854
rect 505102 438618 524546 438854
rect 524782 438618 524866 438854
rect 525102 438618 544546 438854
rect 544782 438618 544866 438854
rect 545102 438618 564546 438854
rect 564782 438618 564866 438854
rect 565102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 826 435454
rect 1062 435218 1146 435454
rect 1382 435218 20826 435454
rect 21062 435218 21146 435454
rect 21382 435218 40826 435454
rect 41062 435218 41146 435454
rect 41382 435218 60826 435454
rect 61062 435218 61146 435454
rect 61382 435218 80826 435454
rect 81062 435218 81146 435454
rect 81382 435218 100826 435454
rect 101062 435218 101146 435454
rect 101382 435218 120826 435454
rect 121062 435218 121146 435454
rect 121382 435218 140826 435454
rect 141062 435218 141146 435454
rect 141382 435218 160826 435454
rect 161062 435218 161146 435454
rect 161382 435218 180826 435454
rect 181062 435218 181146 435454
rect 181382 435218 200826 435454
rect 201062 435218 201146 435454
rect 201382 435218 220826 435454
rect 221062 435218 221146 435454
rect 221382 435218 240826 435454
rect 241062 435218 241146 435454
rect 241382 435218 260826 435454
rect 261062 435218 261146 435454
rect 261382 435218 280826 435454
rect 281062 435218 281146 435454
rect 281382 435218 300826 435454
rect 301062 435218 301146 435454
rect 301382 435218 320826 435454
rect 321062 435218 321146 435454
rect 321382 435218 340826 435454
rect 341062 435218 341146 435454
rect 341382 435218 360826 435454
rect 361062 435218 361146 435454
rect 361382 435218 380826 435454
rect 381062 435218 381146 435454
rect 381382 435218 400826 435454
rect 401062 435218 401146 435454
rect 401382 435218 420826 435454
rect 421062 435218 421146 435454
rect 421382 435218 440826 435454
rect 441062 435218 441146 435454
rect 441382 435218 460826 435454
rect 461062 435218 461146 435454
rect 461382 435218 480826 435454
rect 481062 435218 481146 435454
rect 481382 435218 500826 435454
rect 501062 435218 501146 435454
rect 501382 435218 520826 435454
rect 521062 435218 521146 435454
rect 521382 435218 540826 435454
rect 541062 435218 541146 435454
rect 541382 435218 560826 435454
rect 561062 435218 561146 435454
rect 561382 435218 580826 435454
rect 581062 435218 581146 435454
rect 581382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 826 435134
rect 1062 434898 1146 435134
rect 1382 434898 20826 435134
rect 21062 434898 21146 435134
rect 21382 434898 40826 435134
rect 41062 434898 41146 435134
rect 41382 434898 60826 435134
rect 61062 434898 61146 435134
rect 61382 434898 80826 435134
rect 81062 434898 81146 435134
rect 81382 434898 100826 435134
rect 101062 434898 101146 435134
rect 101382 434898 120826 435134
rect 121062 434898 121146 435134
rect 121382 434898 140826 435134
rect 141062 434898 141146 435134
rect 141382 434898 160826 435134
rect 161062 434898 161146 435134
rect 161382 434898 180826 435134
rect 181062 434898 181146 435134
rect 181382 434898 200826 435134
rect 201062 434898 201146 435134
rect 201382 434898 220826 435134
rect 221062 434898 221146 435134
rect 221382 434898 240826 435134
rect 241062 434898 241146 435134
rect 241382 434898 260826 435134
rect 261062 434898 261146 435134
rect 261382 434898 280826 435134
rect 281062 434898 281146 435134
rect 281382 434898 300826 435134
rect 301062 434898 301146 435134
rect 301382 434898 320826 435134
rect 321062 434898 321146 435134
rect 321382 434898 340826 435134
rect 341062 434898 341146 435134
rect 341382 434898 360826 435134
rect 361062 434898 361146 435134
rect 361382 434898 380826 435134
rect 381062 434898 381146 435134
rect 381382 434898 400826 435134
rect 401062 434898 401146 435134
rect 401382 434898 420826 435134
rect 421062 434898 421146 435134
rect 421382 434898 440826 435134
rect 441062 434898 441146 435134
rect 441382 434898 460826 435134
rect 461062 434898 461146 435134
rect 461382 434898 480826 435134
rect 481062 434898 481146 435134
rect 481382 434898 500826 435134
rect 501062 434898 501146 435134
rect 501382 434898 520826 435134
rect 521062 434898 521146 435134
rect 521382 434898 540826 435134
rect 541062 434898 541146 435134
rect 541382 434898 560826 435134
rect 561062 434898 561146 435134
rect 561382 434898 580826 435134
rect 581062 434898 581146 435134
rect 581382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 21986 428614
rect 22222 428378 22306 428614
rect 22542 428378 41986 428614
rect 42222 428378 42306 428614
rect 42542 428378 61986 428614
rect 62222 428378 62306 428614
rect 62542 428378 81986 428614
rect 82222 428378 82306 428614
rect 82542 428378 101986 428614
rect 102222 428378 102306 428614
rect 102542 428378 121986 428614
rect 122222 428378 122306 428614
rect 122542 428378 141986 428614
rect 142222 428378 142306 428614
rect 142542 428378 161986 428614
rect 162222 428378 162306 428614
rect 162542 428378 181986 428614
rect 182222 428378 182306 428614
rect 182542 428378 201986 428614
rect 202222 428378 202306 428614
rect 202542 428378 221986 428614
rect 222222 428378 222306 428614
rect 222542 428378 241986 428614
rect 242222 428378 242306 428614
rect 242542 428378 261986 428614
rect 262222 428378 262306 428614
rect 262542 428378 281986 428614
rect 282222 428378 282306 428614
rect 282542 428378 301986 428614
rect 302222 428378 302306 428614
rect 302542 428378 321986 428614
rect 322222 428378 322306 428614
rect 322542 428378 341986 428614
rect 342222 428378 342306 428614
rect 342542 428378 361986 428614
rect 362222 428378 362306 428614
rect 362542 428378 381986 428614
rect 382222 428378 382306 428614
rect 382542 428378 401986 428614
rect 402222 428378 402306 428614
rect 402542 428378 421986 428614
rect 422222 428378 422306 428614
rect 422542 428378 441986 428614
rect 442222 428378 442306 428614
rect 442542 428378 461986 428614
rect 462222 428378 462306 428614
rect 462542 428378 481986 428614
rect 482222 428378 482306 428614
rect 482542 428378 501986 428614
rect 502222 428378 502306 428614
rect 502542 428378 521986 428614
rect 522222 428378 522306 428614
rect 522542 428378 541986 428614
rect 542222 428378 542306 428614
rect 542542 428378 561986 428614
rect 562222 428378 562306 428614
rect 562542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 21986 428294
rect 22222 428058 22306 428294
rect 22542 428058 41986 428294
rect 42222 428058 42306 428294
rect 42542 428058 61986 428294
rect 62222 428058 62306 428294
rect 62542 428058 81986 428294
rect 82222 428058 82306 428294
rect 82542 428058 101986 428294
rect 102222 428058 102306 428294
rect 102542 428058 121986 428294
rect 122222 428058 122306 428294
rect 122542 428058 141986 428294
rect 142222 428058 142306 428294
rect 142542 428058 161986 428294
rect 162222 428058 162306 428294
rect 162542 428058 181986 428294
rect 182222 428058 182306 428294
rect 182542 428058 201986 428294
rect 202222 428058 202306 428294
rect 202542 428058 221986 428294
rect 222222 428058 222306 428294
rect 222542 428058 241986 428294
rect 242222 428058 242306 428294
rect 242542 428058 261986 428294
rect 262222 428058 262306 428294
rect 262542 428058 281986 428294
rect 282222 428058 282306 428294
rect 282542 428058 301986 428294
rect 302222 428058 302306 428294
rect 302542 428058 321986 428294
rect 322222 428058 322306 428294
rect 322542 428058 341986 428294
rect 342222 428058 342306 428294
rect 342542 428058 361986 428294
rect 362222 428058 362306 428294
rect 362542 428058 381986 428294
rect 382222 428058 382306 428294
rect 382542 428058 401986 428294
rect 402222 428058 402306 428294
rect 402542 428058 421986 428294
rect 422222 428058 422306 428294
rect 422542 428058 441986 428294
rect 442222 428058 442306 428294
rect 442542 428058 461986 428294
rect 462222 428058 462306 428294
rect 462542 428058 481986 428294
rect 482222 428058 482306 428294
rect 482542 428058 501986 428294
rect 502222 428058 502306 428294
rect 502542 428058 521986 428294
rect 522222 428058 522306 428294
rect 522542 428058 541986 428294
rect 542222 428058 542306 428294
rect 542542 428058 561986 428294
rect 562222 428058 562306 428294
rect 562542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 18266 424894
rect 18502 424658 18586 424894
rect 18822 424658 38266 424894
rect 38502 424658 38586 424894
rect 38822 424658 58266 424894
rect 58502 424658 58586 424894
rect 58822 424658 78266 424894
rect 78502 424658 78586 424894
rect 78822 424658 98266 424894
rect 98502 424658 98586 424894
rect 98822 424658 118266 424894
rect 118502 424658 118586 424894
rect 118822 424658 138266 424894
rect 138502 424658 138586 424894
rect 138822 424658 158266 424894
rect 158502 424658 158586 424894
rect 158822 424658 178266 424894
rect 178502 424658 178586 424894
rect 178822 424658 198266 424894
rect 198502 424658 198586 424894
rect 198822 424658 218266 424894
rect 218502 424658 218586 424894
rect 218822 424658 238266 424894
rect 238502 424658 238586 424894
rect 238822 424658 258266 424894
rect 258502 424658 258586 424894
rect 258822 424658 278266 424894
rect 278502 424658 278586 424894
rect 278822 424658 298266 424894
rect 298502 424658 298586 424894
rect 298822 424658 318266 424894
rect 318502 424658 318586 424894
rect 318822 424658 338266 424894
rect 338502 424658 338586 424894
rect 338822 424658 358266 424894
rect 358502 424658 358586 424894
rect 358822 424658 378266 424894
rect 378502 424658 378586 424894
rect 378822 424658 398266 424894
rect 398502 424658 398586 424894
rect 398822 424658 418266 424894
rect 418502 424658 418586 424894
rect 418822 424658 438266 424894
rect 438502 424658 438586 424894
rect 438822 424658 458266 424894
rect 458502 424658 458586 424894
rect 458822 424658 478266 424894
rect 478502 424658 478586 424894
rect 478822 424658 498266 424894
rect 498502 424658 498586 424894
rect 498822 424658 518266 424894
rect 518502 424658 518586 424894
rect 518822 424658 538266 424894
rect 538502 424658 538586 424894
rect 538822 424658 558266 424894
rect 558502 424658 558586 424894
rect 558822 424658 578266 424894
rect 578502 424658 578586 424894
rect 578822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 18266 424574
rect 18502 424338 18586 424574
rect 18822 424338 38266 424574
rect 38502 424338 38586 424574
rect 38822 424338 58266 424574
rect 58502 424338 58586 424574
rect 58822 424338 78266 424574
rect 78502 424338 78586 424574
rect 78822 424338 98266 424574
rect 98502 424338 98586 424574
rect 98822 424338 118266 424574
rect 118502 424338 118586 424574
rect 118822 424338 138266 424574
rect 138502 424338 138586 424574
rect 138822 424338 158266 424574
rect 158502 424338 158586 424574
rect 158822 424338 178266 424574
rect 178502 424338 178586 424574
rect 178822 424338 198266 424574
rect 198502 424338 198586 424574
rect 198822 424338 218266 424574
rect 218502 424338 218586 424574
rect 218822 424338 238266 424574
rect 238502 424338 238586 424574
rect 238822 424338 258266 424574
rect 258502 424338 258586 424574
rect 258822 424338 278266 424574
rect 278502 424338 278586 424574
rect 278822 424338 298266 424574
rect 298502 424338 298586 424574
rect 298822 424338 318266 424574
rect 318502 424338 318586 424574
rect 318822 424338 338266 424574
rect 338502 424338 338586 424574
rect 338822 424338 358266 424574
rect 358502 424338 358586 424574
rect 358822 424338 378266 424574
rect 378502 424338 378586 424574
rect 378822 424338 398266 424574
rect 398502 424338 398586 424574
rect 398822 424338 418266 424574
rect 418502 424338 418586 424574
rect 418822 424338 438266 424574
rect 438502 424338 438586 424574
rect 438822 424338 458266 424574
rect 458502 424338 458586 424574
rect 458822 424338 478266 424574
rect 478502 424338 478586 424574
rect 478822 424338 498266 424574
rect 498502 424338 498586 424574
rect 498822 424338 518266 424574
rect 518502 424338 518586 424574
rect 518822 424338 538266 424574
rect 538502 424338 538586 424574
rect 538822 424338 558266 424574
rect 558502 424338 558586 424574
rect 558822 424338 578266 424574
rect 578502 424338 578586 424574
rect 578822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 14546 421174
rect 14782 420938 14866 421174
rect 15102 420938 34546 421174
rect 34782 420938 34866 421174
rect 35102 420938 54546 421174
rect 54782 420938 54866 421174
rect 55102 420938 74546 421174
rect 74782 420938 74866 421174
rect 75102 420938 94546 421174
rect 94782 420938 94866 421174
rect 95102 420938 114546 421174
rect 114782 420938 114866 421174
rect 115102 420938 134546 421174
rect 134782 420938 134866 421174
rect 135102 420938 154546 421174
rect 154782 420938 154866 421174
rect 155102 420938 174546 421174
rect 174782 420938 174866 421174
rect 175102 420938 194546 421174
rect 194782 420938 194866 421174
rect 195102 420938 214546 421174
rect 214782 420938 214866 421174
rect 215102 420938 234546 421174
rect 234782 420938 234866 421174
rect 235102 420938 254546 421174
rect 254782 420938 254866 421174
rect 255102 420938 274546 421174
rect 274782 420938 274866 421174
rect 275102 420938 294546 421174
rect 294782 420938 294866 421174
rect 295102 420938 314546 421174
rect 314782 420938 314866 421174
rect 315102 420938 334546 421174
rect 334782 420938 334866 421174
rect 335102 420938 354546 421174
rect 354782 420938 354866 421174
rect 355102 420938 374546 421174
rect 374782 420938 374866 421174
rect 375102 420938 394546 421174
rect 394782 420938 394866 421174
rect 395102 420938 414546 421174
rect 414782 420938 414866 421174
rect 415102 420938 434546 421174
rect 434782 420938 434866 421174
rect 435102 420938 454546 421174
rect 454782 420938 454866 421174
rect 455102 420938 474546 421174
rect 474782 420938 474866 421174
rect 475102 420938 494546 421174
rect 494782 420938 494866 421174
rect 495102 420938 514546 421174
rect 514782 420938 514866 421174
rect 515102 420938 534546 421174
rect 534782 420938 534866 421174
rect 535102 420938 554546 421174
rect 554782 420938 554866 421174
rect 555102 420938 574546 421174
rect 574782 420938 574866 421174
rect 575102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 14546 420854
rect 14782 420618 14866 420854
rect 15102 420618 34546 420854
rect 34782 420618 34866 420854
rect 35102 420618 54546 420854
rect 54782 420618 54866 420854
rect 55102 420618 74546 420854
rect 74782 420618 74866 420854
rect 75102 420618 94546 420854
rect 94782 420618 94866 420854
rect 95102 420618 114546 420854
rect 114782 420618 114866 420854
rect 115102 420618 134546 420854
rect 134782 420618 134866 420854
rect 135102 420618 154546 420854
rect 154782 420618 154866 420854
rect 155102 420618 174546 420854
rect 174782 420618 174866 420854
rect 175102 420618 194546 420854
rect 194782 420618 194866 420854
rect 195102 420618 214546 420854
rect 214782 420618 214866 420854
rect 215102 420618 234546 420854
rect 234782 420618 234866 420854
rect 235102 420618 254546 420854
rect 254782 420618 254866 420854
rect 255102 420618 274546 420854
rect 274782 420618 274866 420854
rect 275102 420618 294546 420854
rect 294782 420618 294866 420854
rect 295102 420618 314546 420854
rect 314782 420618 314866 420854
rect 315102 420618 334546 420854
rect 334782 420618 334866 420854
rect 335102 420618 354546 420854
rect 354782 420618 354866 420854
rect 355102 420618 374546 420854
rect 374782 420618 374866 420854
rect 375102 420618 394546 420854
rect 394782 420618 394866 420854
rect 395102 420618 414546 420854
rect 414782 420618 414866 420854
rect 415102 420618 434546 420854
rect 434782 420618 434866 420854
rect 435102 420618 454546 420854
rect 454782 420618 454866 420854
rect 455102 420618 474546 420854
rect 474782 420618 474866 420854
rect 475102 420618 494546 420854
rect 494782 420618 494866 420854
rect 495102 420618 514546 420854
rect 514782 420618 514866 420854
rect 515102 420618 534546 420854
rect 534782 420618 534866 420854
rect 535102 420618 554546 420854
rect 554782 420618 554866 420854
rect 555102 420618 574546 420854
rect 574782 420618 574866 420854
rect 575102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 10826 417454
rect 11062 417218 11146 417454
rect 11382 417218 30826 417454
rect 31062 417218 31146 417454
rect 31382 417218 50826 417454
rect 51062 417218 51146 417454
rect 51382 417218 70826 417454
rect 71062 417218 71146 417454
rect 71382 417218 90826 417454
rect 91062 417218 91146 417454
rect 91382 417218 110826 417454
rect 111062 417218 111146 417454
rect 111382 417218 130826 417454
rect 131062 417218 131146 417454
rect 131382 417218 150826 417454
rect 151062 417218 151146 417454
rect 151382 417218 170826 417454
rect 171062 417218 171146 417454
rect 171382 417218 190826 417454
rect 191062 417218 191146 417454
rect 191382 417218 210826 417454
rect 211062 417218 211146 417454
rect 211382 417218 230826 417454
rect 231062 417218 231146 417454
rect 231382 417218 250826 417454
rect 251062 417218 251146 417454
rect 251382 417218 270826 417454
rect 271062 417218 271146 417454
rect 271382 417218 290826 417454
rect 291062 417218 291146 417454
rect 291382 417218 310826 417454
rect 311062 417218 311146 417454
rect 311382 417218 330826 417454
rect 331062 417218 331146 417454
rect 331382 417218 350826 417454
rect 351062 417218 351146 417454
rect 351382 417218 370826 417454
rect 371062 417218 371146 417454
rect 371382 417218 390826 417454
rect 391062 417218 391146 417454
rect 391382 417218 410826 417454
rect 411062 417218 411146 417454
rect 411382 417218 430826 417454
rect 431062 417218 431146 417454
rect 431382 417218 450826 417454
rect 451062 417218 451146 417454
rect 451382 417218 470826 417454
rect 471062 417218 471146 417454
rect 471382 417218 490826 417454
rect 491062 417218 491146 417454
rect 491382 417218 510826 417454
rect 511062 417218 511146 417454
rect 511382 417218 530826 417454
rect 531062 417218 531146 417454
rect 531382 417218 550826 417454
rect 551062 417218 551146 417454
rect 551382 417218 570826 417454
rect 571062 417218 571146 417454
rect 571382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 10826 417134
rect 11062 416898 11146 417134
rect 11382 416898 30826 417134
rect 31062 416898 31146 417134
rect 31382 416898 50826 417134
rect 51062 416898 51146 417134
rect 51382 416898 70826 417134
rect 71062 416898 71146 417134
rect 71382 416898 90826 417134
rect 91062 416898 91146 417134
rect 91382 416898 110826 417134
rect 111062 416898 111146 417134
rect 111382 416898 130826 417134
rect 131062 416898 131146 417134
rect 131382 416898 150826 417134
rect 151062 416898 151146 417134
rect 151382 416898 170826 417134
rect 171062 416898 171146 417134
rect 171382 416898 190826 417134
rect 191062 416898 191146 417134
rect 191382 416898 210826 417134
rect 211062 416898 211146 417134
rect 211382 416898 230826 417134
rect 231062 416898 231146 417134
rect 231382 416898 250826 417134
rect 251062 416898 251146 417134
rect 251382 416898 270826 417134
rect 271062 416898 271146 417134
rect 271382 416898 290826 417134
rect 291062 416898 291146 417134
rect 291382 416898 310826 417134
rect 311062 416898 311146 417134
rect 311382 416898 330826 417134
rect 331062 416898 331146 417134
rect 331382 416898 350826 417134
rect 351062 416898 351146 417134
rect 351382 416898 370826 417134
rect 371062 416898 371146 417134
rect 371382 416898 390826 417134
rect 391062 416898 391146 417134
rect 391382 416898 410826 417134
rect 411062 416898 411146 417134
rect 411382 416898 430826 417134
rect 431062 416898 431146 417134
rect 431382 416898 450826 417134
rect 451062 416898 451146 417134
rect 451382 416898 470826 417134
rect 471062 416898 471146 417134
rect 471382 416898 490826 417134
rect 491062 416898 491146 417134
rect 491382 416898 510826 417134
rect 511062 416898 511146 417134
rect 511382 416898 530826 417134
rect 531062 416898 531146 417134
rect 531382 416898 550826 417134
rect 551062 416898 551146 417134
rect 551382 416898 570826 417134
rect 571062 416898 571146 417134
rect 571382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 11986 410614
rect 12222 410378 12306 410614
rect 12542 410378 31986 410614
rect 32222 410378 32306 410614
rect 32542 410378 51986 410614
rect 52222 410378 52306 410614
rect 52542 410378 71986 410614
rect 72222 410378 72306 410614
rect 72542 410378 91986 410614
rect 92222 410378 92306 410614
rect 92542 410378 111986 410614
rect 112222 410378 112306 410614
rect 112542 410378 131986 410614
rect 132222 410378 132306 410614
rect 132542 410378 151986 410614
rect 152222 410378 152306 410614
rect 152542 410378 171986 410614
rect 172222 410378 172306 410614
rect 172542 410378 191986 410614
rect 192222 410378 192306 410614
rect 192542 410378 211986 410614
rect 212222 410378 212306 410614
rect 212542 410378 231986 410614
rect 232222 410378 232306 410614
rect 232542 410378 251986 410614
rect 252222 410378 252306 410614
rect 252542 410378 271986 410614
rect 272222 410378 272306 410614
rect 272542 410378 291986 410614
rect 292222 410378 292306 410614
rect 292542 410378 311986 410614
rect 312222 410378 312306 410614
rect 312542 410378 331986 410614
rect 332222 410378 332306 410614
rect 332542 410378 351986 410614
rect 352222 410378 352306 410614
rect 352542 410378 371986 410614
rect 372222 410378 372306 410614
rect 372542 410378 391986 410614
rect 392222 410378 392306 410614
rect 392542 410378 411986 410614
rect 412222 410378 412306 410614
rect 412542 410378 431986 410614
rect 432222 410378 432306 410614
rect 432542 410378 451986 410614
rect 452222 410378 452306 410614
rect 452542 410378 471986 410614
rect 472222 410378 472306 410614
rect 472542 410378 491986 410614
rect 492222 410378 492306 410614
rect 492542 410378 511986 410614
rect 512222 410378 512306 410614
rect 512542 410378 531986 410614
rect 532222 410378 532306 410614
rect 532542 410378 551986 410614
rect 552222 410378 552306 410614
rect 552542 410378 571986 410614
rect 572222 410378 572306 410614
rect 572542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 11986 410294
rect 12222 410058 12306 410294
rect 12542 410058 31986 410294
rect 32222 410058 32306 410294
rect 32542 410058 51986 410294
rect 52222 410058 52306 410294
rect 52542 410058 71986 410294
rect 72222 410058 72306 410294
rect 72542 410058 91986 410294
rect 92222 410058 92306 410294
rect 92542 410058 111986 410294
rect 112222 410058 112306 410294
rect 112542 410058 131986 410294
rect 132222 410058 132306 410294
rect 132542 410058 151986 410294
rect 152222 410058 152306 410294
rect 152542 410058 171986 410294
rect 172222 410058 172306 410294
rect 172542 410058 191986 410294
rect 192222 410058 192306 410294
rect 192542 410058 211986 410294
rect 212222 410058 212306 410294
rect 212542 410058 231986 410294
rect 232222 410058 232306 410294
rect 232542 410058 251986 410294
rect 252222 410058 252306 410294
rect 252542 410058 271986 410294
rect 272222 410058 272306 410294
rect 272542 410058 291986 410294
rect 292222 410058 292306 410294
rect 292542 410058 311986 410294
rect 312222 410058 312306 410294
rect 312542 410058 331986 410294
rect 332222 410058 332306 410294
rect 332542 410058 351986 410294
rect 352222 410058 352306 410294
rect 352542 410058 371986 410294
rect 372222 410058 372306 410294
rect 372542 410058 391986 410294
rect 392222 410058 392306 410294
rect 392542 410058 411986 410294
rect 412222 410058 412306 410294
rect 412542 410058 431986 410294
rect 432222 410058 432306 410294
rect 432542 410058 451986 410294
rect 452222 410058 452306 410294
rect 452542 410058 471986 410294
rect 472222 410058 472306 410294
rect 472542 410058 491986 410294
rect 492222 410058 492306 410294
rect 492542 410058 511986 410294
rect 512222 410058 512306 410294
rect 512542 410058 531986 410294
rect 532222 410058 532306 410294
rect 532542 410058 551986 410294
rect 552222 410058 552306 410294
rect 552542 410058 571986 410294
rect 572222 410058 572306 410294
rect 572542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 8266 406894
rect 8502 406658 8586 406894
rect 8822 406658 28266 406894
rect 28502 406658 28586 406894
rect 28822 406658 48266 406894
rect 48502 406658 48586 406894
rect 48822 406658 68266 406894
rect 68502 406658 68586 406894
rect 68822 406658 88266 406894
rect 88502 406658 88586 406894
rect 88822 406658 108266 406894
rect 108502 406658 108586 406894
rect 108822 406658 128266 406894
rect 128502 406658 128586 406894
rect 128822 406658 148266 406894
rect 148502 406658 148586 406894
rect 148822 406658 168266 406894
rect 168502 406658 168586 406894
rect 168822 406658 188266 406894
rect 188502 406658 188586 406894
rect 188822 406658 208266 406894
rect 208502 406658 208586 406894
rect 208822 406658 228266 406894
rect 228502 406658 228586 406894
rect 228822 406658 248266 406894
rect 248502 406658 248586 406894
rect 248822 406658 268266 406894
rect 268502 406658 268586 406894
rect 268822 406658 288266 406894
rect 288502 406658 288586 406894
rect 288822 406658 308266 406894
rect 308502 406658 308586 406894
rect 308822 406658 328266 406894
rect 328502 406658 328586 406894
rect 328822 406658 348266 406894
rect 348502 406658 348586 406894
rect 348822 406658 368266 406894
rect 368502 406658 368586 406894
rect 368822 406658 388266 406894
rect 388502 406658 388586 406894
rect 388822 406658 408266 406894
rect 408502 406658 408586 406894
rect 408822 406658 428266 406894
rect 428502 406658 428586 406894
rect 428822 406658 448266 406894
rect 448502 406658 448586 406894
rect 448822 406658 468266 406894
rect 468502 406658 468586 406894
rect 468822 406658 488266 406894
rect 488502 406658 488586 406894
rect 488822 406658 508266 406894
rect 508502 406658 508586 406894
rect 508822 406658 528266 406894
rect 528502 406658 528586 406894
rect 528822 406658 548266 406894
rect 548502 406658 548586 406894
rect 548822 406658 568266 406894
rect 568502 406658 568586 406894
rect 568822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 8266 406574
rect 8502 406338 8586 406574
rect 8822 406338 28266 406574
rect 28502 406338 28586 406574
rect 28822 406338 48266 406574
rect 48502 406338 48586 406574
rect 48822 406338 68266 406574
rect 68502 406338 68586 406574
rect 68822 406338 88266 406574
rect 88502 406338 88586 406574
rect 88822 406338 108266 406574
rect 108502 406338 108586 406574
rect 108822 406338 128266 406574
rect 128502 406338 128586 406574
rect 128822 406338 148266 406574
rect 148502 406338 148586 406574
rect 148822 406338 168266 406574
rect 168502 406338 168586 406574
rect 168822 406338 188266 406574
rect 188502 406338 188586 406574
rect 188822 406338 208266 406574
rect 208502 406338 208586 406574
rect 208822 406338 228266 406574
rect 228502 406338 228586 406574
rect 228822 406338 248266 406574
rect 248502 406338 248586 406574
rect 248822 406338 268266 406574
rect 268502 406338 268586 406574
rect 268822 406338 288266 406574
rect 288502 406338 288586 406574
rect 288822 406338 308266 406574
rect 308502 406338 308586 406574
rect 308822 406338 328266 406574
rect 328502 406338 328586 406574
rect 328822 406338 348266 406574
rect 348502 406338 348586 406574
rect 348822 406338 368266 406574
rect 368502 406338 368586 406574
rect 368822 406338 388266 406574
rect 388502 406338 388586 406574
rect 388822 406338 408266 406574
rect 408502 406338 408586 406574
rect 408822 406338 428266 406574
rect 428502 406338 428586 406574
rect 428822 406338 448266 406574
rect 448502 406338 448586 406574
rect 448822 406338 468266 406574
rect 468502 406338 468586 406574
rect 468822 406338 488266 406574
rect 488502 406338 488586 406574
rect 488822 406338 508266 406574
rect 508502 406338 508586 406574
rect 508822 406338 528266 406574
rect 528502 406338 528586 406574
rect 528822 406338 548266 406574
rect 548502 406338 548586 406574
rect 548822 406338 568266 406574
rect 568502 406338 568586 406574
rect 568822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 4546 403174
rect 4782 402938 4866 403174
rect 5102 402938 24546 403174
rect 24782 402938 24866 403174
rect 25102 402938 44546 403174
rect 44782 402938 44866 403174
rect 45102 402938 64546 403174
rect 64782 402938 64866 403174
rect 65102 402938 84546 403174
rect 84782 402938 84866 403174
rect 85102 402938 104546 403174
rect 104782 402938 104866 403174
rect 105102 402938 124546 403174
rect 124782 402938 124866 403174
rect 125102 402938 144546 403174
rect 144782 402938 144866 403174
rect 145102 402938 164546 403174
rect 164782 402938 164866 403174
rect 165102 402938 184546 403174
rect 184782 402938 184866 403174
rect 185102 402938 204546 403174
rect 204782 402938 204866 403174
rect 205102 402938 224546 403174
rect 224782 402938 224866 403174
rect 225102 402938 244546 403174
rect 244782 402938 244866 403174
rect 245102 402938 264546 403174
rect 264782 402938 264866 403174
rect 265102 402938 284546 403174
rect 284782 402938 284866 403174
rect 285102 402938 304546 403174
rect 304782 402938 304866 403174
rect 305102 402938 324546 403174
rect 324782 402938 324866 403174
rect 325102 402938 344546 403174
rect 344782 402938 344866 403174
rect 345102 402938 364546 403174
rect 364782 402938 364866 403174
rect 365102 402938 384546 403174
rect 384782 402938 384866 403174
rect 385102 402938 404546 403174
rect 404782 402938 404866 403174
rect 405102 402938 424546 403174
rect 424782 402938 424866 403174
rect 425102 402938 444546 403174
rect 444782 402938 444866 403174
rect 445102 402938 464546 403174
rect 464782 402938 464866 403174
rect 465102 402938 484546 403174
rect 484782 402938 484866 403174
rect 485102 402938 504546 403174
rect 504782 402938 504866 403174
rect 505102 402938 524546 403174
rect 524782 402938 524866 403174
rect 525102 402938 544546 403174
rect 544782 402938 544866 403174
rect 545102 402938 564546 403174
rect 564782 402938 564866 403174
rect 565102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 4546 402854
rect 4782 402618 4866 402854
rect 5102 402618 24546 402854
rect 24782 402618 24866 402854
rect 25102 402618 44546 402854
rect 44782 402618 44866 402854
rect 45102 402618 64546 402854
rect 64782 402618 64866 402854
rect 65102 402618 84546 402854
rect 84782 402618 84866 402854
rect 85102 402618 104546 402854
rect 104782 402618 104866 402854
rect 105102 402618 124546 402854
rect 124782 402618 124866 402854
rect 125102 402618 144546 402854
rect 144782 402618 144866 402854
rect 145102 402618 164546 402854
rect 164782 402618 164866 402854
rect 165102 402618 184546 402854
rect 184782 402618 184866 402854
rect 185102 402618 204546 402854
rect 204782 402618 204866 402854
rect 205102 402618 224546 402854
rect 224782 402618 224866 402854
rect 225102 402618 244546 402854
rect 244782 402618 244866 402854
rect 245102 402618 264546 402854
rect 264782 402618 264866 402854
rect 265102 402618 284546 402854
rect 284782 402618 284866 402854
rect 285102 402618 304546 402854
rect 304782 402618 304866 402854
rect 305102 402618 324546 402854
rect 324782 402618 324866 402854
rect 325102 402618 344546 402854
rect 344782 402618 344866 402854
rect 345102 402618 364546 402854
rect 364782 402618 364866 402854
rect 365102 402618 384546 402854
rect 384782 402618 384866 402854
rect 385102 402618 404546 402854
rect 404782 402618 404866 402854
rect 405102 402618 424546 402854
rect 424782 402618 424866 402854
rect 425102 402618 444546 402854
rect 444782 402618 444866 402854
rect 445102 402618 464546 402854
rect 464782 402618 464866 402854
rect 465102 402618 484546 402854
rect 484782 402618 484866 402854
rect 485102 402618 504546 402854
rect 504782 402618 504866 402854
rect 505102 402618 524546 402854
rect 524782 402618 524866 402854
rect 525102 402618 544546 402854
rect 544782 402618 544866 402854
rect 545102 402618 564546 402854
rect 564782 402618 564866 402854
rect 565102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 826 399454
rect 1062 399218 1146 399454
rect 1382 399218 20826 399454
rect 21062 399218 21146 399454
rect 21382 399218 40826 399454
rect 41062 399218 41146 399454
rect 41382 399218 60826 399454
rect 61062 399218 61146 399454
rect 61382 399218 80826 399454
rect 81062 399218 81146 399454
rect 81382 399218 100826 399454
rect 101062 399218 101146 399454
rect 101382 399218 120826 399454
rect 121062 399218 121146 399454
rect 121382 399218 140826 399454
rect 141062 399218 141146 399454
rect 141382 399218 160826 399454
rect 161062 399218 161146 399454
rect 161382 399218 180826 399454
rect 181062 399218 181146 399454
rect 181382 399218 200826 399454
rect 201062 399218 201146 399454
rect 201382 399218 220826 399454
rect 221062 399218 221146 399454
rect 221382 399218 240826 399454
rect 241062 399218 241146 399454
rect 241382 399218 260826 399454
rect 261062 399218 261146 399454
rect 261382 399218 280826 399454
rect 281062 399218 281146 399454
rect 281382 399218 300826 399454
rect 301062 399218 301146 399454
rect 301382 399218 320826 399454
rect 321062 399218 321146 399454
rect 321382 399218 340826 399454
rect 341062 399218 341146 399454
rect 341382 399218 360826 399454
rect 361062 399218 361146 399454
rect 361382 399218 380826 399454
rect 381062 399218 381146 399454
rect 381382 399218 400826 399454
rect 401062 399218 401146 399454
rect 401382 399218 420826 399454
rect 421062 399218 421146 399454
rect 421382 399218 440826 399454
rect 441062 399218 441146 399454
rect 441382 399218 460826 399454
rect 461062 399218 461146 399454
rect 461382 399218 480826 399454
rect 481062 399218 481146 399454
rect 481382 399218 500826 399454
rect 501062 399218 501146 399454
rect 501382 399218 520826 399454
rect 521062 399218 521146 399454
rect 521382 399218 540826 399454
rect 541062 399218 541146 399454
rect 541382 399218 560826 399454
rect 561062 399218 561146 399454
rect 561382 399218 580826 399454
rect 581062 399218 581146 399454
rect 581382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 826 399134
rect 1062 398898 1146 399134
rect 1382 398898 20826 399134
rect 21062 398898 21146 399134
rect 21382 398898 40826 399134
rect 41062 398898 41146 399134
rect 41382 398898 60826 399134
rect 61062 398898 61146 399134
rect 61382 398898 80826 399134
rect 81062 398898 81146 399134
rect 81382 398898 100826 399134
rect 101062 398898 101146 399134
rect 101382 398898 120826 399134
rect 121062 398898 121146 399134
rect 121382 398898 140826 399134
rect 141062 398898 141146 399134
rect 141382 398898 160826 399134
rect 161062 398898 161146 399134
rect 161382 398898 180826 399134
rect 181062 398898 181146 399134
rect 181382 398898 200826 399134
rect 201062 398898 201146 399134
rect 201382 398898 220826 399134
rect 221062 398898 221146 399134
rect 221382 398898 240826 399134
rect 241062 398898 241146 399134
rect 241382 398898 260826 399134
rect 261062 398898 261146 399134
rect 261382 398898 280826 399134
rect 281062 398898 281146 399134
rect 281382 398898 300826 399134
rect 301062 398898 301146 399134
rect 301382 398898 320826 399134
rect 321062 398898 321146 399134
rect 321382 398898 340826 399134
rect 341062 398898 341146 399134
rect 341382 398898 360826 399134
rect 361062 398898 361146 399134
rect 361382 398898 380826 399134
rect 381062 398898 381146 399134
rect 381382 398898 400826 399134
rect 401062 398898 401146 399134
rect 401382 398898 420826 399134
rect 421062 398898 421146 399134
rect 421382 398898 440826 399134
rect 441062 398898 441146 399134
rect 441382 398898 460826 399134
rect 461062 398898 461146 399134
rect 461382 398898 480826 399134
rect 481062 398898 481146 399134
rect 481382 398898 500826 399134
rect 501062 398898 501146 399134
rect 501382 398898 520826 399134
rect 521062 398898 521146 399134
rect 521382 398898 540826 399134
rect 541062 398898 541146 399134
rect 541382 398898 560826 399134
rect 561062 398898 561146 399134
rect 561382 398898 580826 399134
rect 581062 398898 581146 399134
rect 581382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 21986 392614
rect 22222 392378 22306 392614
rect 22542 392378 41986 392614
rect 42222 392378 42306 392614
rect 42542 392378 61986 392614
rect 62222 392378 62306 392614
rect 62542 392378 81986 392614
rect 82222 392378 82306 392614
rect 82542 392378 101986 392614
rect 102222 392378 102306 392614
rect 102542 392378 121986 392614
rect 122222 392378 122306 392614
rect 122542 392378 141986 392614
rect 142222 392378 142306 392614
rect 142542 392378 161986 392614
rect 162222 392378 162306 392614
rect 162542 392378 181986 392614
rect 182222 392378 182306 392614
rect 182542 392378 201986 392614
rect 202222 392378 202306 392614
rect 202542 392378 221986 392614
rect 222222 392378 222306 392614
rect 222542 392378 241986 392614
rect 242222 392378 242306 392614
rect 242542 392378 261986 392614
rect 262222 392378 262306 392614
rect 262542 392378 281986 392614
rect 282222 392378 282306 392614
rect 282542 392378 301986 392614
rect 302222 392378 302306 392614
rect 302542 392378 321986 392614
rect 322222 392378 322306 392614
rect 322542 392378 341986 392614
rect 342222 392378 342306 392614
rect 342542 392378 361986 392614
rect 362222 392378 362306 392614
rect 362542 392378 381986 392614
rect 382222 392378 382306 392614
rect 382542 392378 401986 392614
rect 402222 392378 402306 392614
rect 402542 392378 421986 392614
rect 422222 392378 422306 392614
rect 422542 392378 441986 392614
rect 442222 392378 442306 392614
rect 442542 392378 461986 392614
rect 462222 392378 462306 392614
rect 462542 392378 481986 392614
rect 482222 392378 482306 392614
rect 482542 392378 501986 392614
rect 502222 392378 502306 392614
rect 502542 392378 521986 392614
rect 522222 392378 522306 392614
rect 522542 392378 541986 392614
rect 542222 392378 542306 392614
rect 542542 392378 561986 392614
rect 562222 392378 562306 392614
rect 562542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 21986 392294
rect 22222 392058 22306 392294
rect 22542 392058 41986 392294
rect 42222 392058 42306 392294
rect 42542 392058 61986 392294
rect 62222 392058 62306 392294
rect 62542 392058 81986 392294
rect 82222 392058 82306 392294
rect 82542 392058 101986 392294
rect 102222 392058 102306 392294
rect 102542 392058 121986 392294
rect 122222 392058 122306 392294
rect 122542 392058 141986 392294
rect 142222 392058 142306 392294
rect 142542 392058 161986 392294
rect 162222 392058 162306 392294
rect 162542 392058 181986 392294
rect 182222 392058 182306 392294
rect 182542 392058 201986 392294
rect 202222 392058 202306 392294
rect 202542 392058 221986 392294
rect 222222 392058 222306 392294
rect 222542 392058 241986 392294
rect 242222 392058 242306 392294
rect 242542 392058 261986 392294
rect 262222 392058 262306 392294
rect 262542 392058 281986 392294
rect 282222 392058 282306 392294
rect 282542 392058 301986 392294
rect 302222 392058 302306 392294
rect 302542 392058 321986 392294
rect 322222 392058 322306 392294
rect 322542 392058 341986 392294
rect 342222 392058 342306 392294
rect 342542 392058 361986 392294
rect 362222 392058 362306 392294
rect 362542 392058 381986 392294
rect 382222 392058 382306 392294
rect 382542 392058 401986 392294
rect 402222 392058 402306 392294
rect 402542 392058 421986 392294
rect 422222 392058 422306 392294
rect 422542 392058 441986 392294
rect 442222 392058 442306 392294
rect 442542 392058 461986 392294
rect 462222 392058 462306 392294
rect 462542 392058 481986 392294
rect 482222 392058 482306 392294
rect 482542 392058 501986 392294
rect 502222 392058 502306 392294
rect 502542 392058 521986 392294
rect 522222 392058 522306 392294
rect 522542 392058 541986 392294
rect 542222 392058 542306 392294
rect 542542 392058 561986 392294
rect 562222 392058 562306 392294
rect 562542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 18266 388894
rect 18502 388658 18586 388894
rect 18822 388658 38266 388894
rect 38502 388658 38586 388894
rect 38822 388658 58266 388894
rect 58502 388658 58586 388894
rect 58822 388658 78266 388894
rect 78502 388658 78586 388894
rect 78822 388658 98266 388894
rect 98502 388658 98586 388894
rect 98822 388658 118266 388894
rect 118502 388658 118586 388894
rect 118822 388658 138266 388894
rect 138502 388658 138586 388894
rect 138822 388658 158266 388894
rect 158502 388658 158586 388894
rect 158822 388658 178266 388894
rect 178502 388658 178586 388894
rect 178822 388658 198266 388894
rect 198502 388658 198586 388894
rect 198822 388658 218266 388894
rect 218502 388658 218586 388894
rect 218822 388658 238266 388894
rect 238502 388658 238586 388894
rect 238822 388658 258266 388894
rect 258502 388658 258586 388894
rect 258822 388658 278266 388894
rect 278502 388658 278586 388894
rect 278822 388658 298266 388894
rect 298502 388658 298586 388894
rect 298822 388658 318266 388894
rect 318502 388658 318586 388894
rect 318822 388658 338266 388894
rect 338502 388658 338586 388894
rect 338822 388658 358266 388894
rect 358502 388658 358586 388894
rect 358822 388658 378266 388894
rect 378502 388658 378586 388894
rect 378822 388658 398266 388894
rect 398502 388658 398586 388894
rect 398822 388658 418266 388894
rect 418502 388658 418586 388894
rect 418822 388658 438266 388894
rect 438502 388658 438586 388894
rect 438822 388658 458266 388894
rect 458502 388658 458586 388894
rect 458822 388658 478266 388894
rect 478502 388658 478586 388894
rect 478822 388658 498266 388894
rect 498502 388658 498586 388894
rect 498822 388658 518266 388894
rect 518502 388658 518586 388894
rect 518822 388658 538266 388894
rect 538502 388658 538586 388894
rect 538822 388658 558266 388894
rect 558502 388658 558586 388894
rect 558822 388658 578266 388894
rect 578502 388658 578586 388894
rect 578822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 18266 388574
rect 18502 388338 18586 388574
rect 18822 388338 38266 388574
rect 38502 388338 38586 388574
rect 38822 388338 58266 388574
rect 58502 388338 58586 388574
rect 58822 388338 78266 388574
rect 78502 388338 78586 388574
rect 78822 388338 98266 388574
rect 98502 388338 98586 388574
rect 98822 388338 118266 388574
rect 118502 388338 118586 388574
rect 118822 388338 138266 388574
rect 138502 388338 138586 388574
rect 138822 388338 158266 388574
rect 158502 388338 158586 388574
rect 158822 388338 178266 388574
rect 178502 388338 178586 388574
rect 178822 388338 198266 388574
rect 198502 388338 198586 388574
rect 198822 388338 218266 388574
rect 218502 388338 218586 388574
rect 218822 388338 238266 388574
rect 238502 388338 238586 388574
rect 238822 388338 258266 388574
rect 258502 388338 258586 388574
rect 258822 388338 278266 388574
rect 278502 388338 278586 388574
rect 278822 388338 298266 388574
rect 298502 388338 298586 388574
rect 298822 388338 318266 388574
rect 318502 388338 318586 388574
rect 318822 388338 338266 388574
rect 338502 388338 338586 388574
rect 338822 388338 358266 388574
rect 358502 388338 358586 388574
rect 358822 388338 378266 388574
rect 378502 388338 378586 388574
rect 378822 388338 398266 388574
rect 398502 388338 398586 388574
rect 398822 388338 418266 388574
rect 418502 388338 418586 388574
rect 418822 388338 438266 388574
rect 438502 388338 438586 388574
rect 438822 388338 458266 388574
rect 458502 388338 458586 388574
rect 458822 388338 478266 388574
rect 478502 388338 478586 388574
rect 478822 388338 498266 388574
rect 498502 388338 498586 388574
rect 498822 388338 518266 388574
rect 518502 388338 518586 388574
rect 518822 388338 538266 388574
rect 538502 388338 538586 388574
rect 538822 388338 558266 388574
rect 558502 388338 558586 388574
rect 558822 388338 578266 388574
rect 578502 388338 578586 388574
rect 578822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 14546 385174
rect 14782 384938 14866 385174
rect 15102 384938 34546 385174
rect 34782 384938 34866 385174
rect 35102 384938 54546 385174
rect 54782 384938 54866 385174
rect 55102 384938 74546 385174
rect 74782 384938 74866 385174
rect 75102 384938 94546 385174
rect 94782 384938 94866 385174
rect 95102 384938 114546 385174
rect 114782 384938 114866 385174
rect 115102 384938 134546 385174
rect 134782 384938 134866 385174
rect 135102 384938 154546 385174
rect 154782 384938 154866 385174
rect 155102 384938 174546 385174
rect 174782 384938 174866 385174
rect 175102 384938 194546 385174
rect 194782 384938 194866 385174
rect 195102 384938 214546 385174
rect 214782 384938 214866 385174
rect 215102 384938 234546 385174
rect 234782 384938 234866 385174
rect 235102 384938 254546 385174
rect 254782 384938 254866 385174
rect 255102 384938 274546 385174
rect 274782 384938 274866 385174
rect 275102 384938 294546 385174
rect 294782 384938 294866 385174
rect 295102 384938 314546 385174
rect 314782 384938 314866 385174
rect 315102 384938 334546 385174
rect 334782 384938 334866 385174
rect 335102 384938 354546 385174
rect 354782 384938 354866 385174
rect 355102 384938 374546 385174
rect 374782 384938 374866 385174
rect 375102 384938 394546 385174
rect 394782 384938 394866 385174
rect 395102 384938 414546 385174
rect 414782 384938 414866 385174
rect 415102 384938 434546 385174
rect 434782 384938 434866 385174
rect 435102 384938 454546 385174
rect 454782 384938 454866 385174
rect 455102 384938 474546 385174
rect 474782 384938 474866 385174
rect 475102 384938 494546 385174
rect 494782 384938 494866 385174
rect 495102 384938 514546 385174
rect 514782 384938 514866 385174
rect 515102 384938 534546 385174
rect 534782 384938 534866 385174
rect 535102 384938 554546 385174
rect 554782 384938 554866 385174
rect 555102 384938 574546 385174
rect 574782 384938 574866 385174
rect 575102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 14546 384854
rect 14782 384618 14866 384854
rect 15102 384618 34546 384854
rect 34782 384618 34866 384854
rect 35102 384618 54546 384854
rect 54782 384618 54866 384854
rect 55102 384618 74546 384854
rect 74782 384618 74866 384854
rect 75102 384618 94546 384854
rect 94782 384618 94866 384854
rect 95102 384618 114546 384854
rect 114782 384618 114866 384854
rect 115102 384618 134546 384854
rect 134782 384618 134866 384854
rect 135102 384618 154546 384854
rect 154782 384618 154866 384854
rect 155102 384618 174546 384854
rect 174782 384618 174866 384854
rect 175102 384618 194546 384854
rect 194782 384618 194866 384854
rect 195102 384618 214546 384854
rect 214782 384618 214866 384854
rect 215102 384618 234546 384854
rect 234782 384618 234866 384854
rect 235102 384618 254546 384854
rect 254782 384618 254866 384854
rect 255102 384618 274546 384854
rect 274782 384618 274866 384854
rect 275102 384618 294546 384854
rect 294782 384618 294866 384854
rect 295102 384618 314546 384854
rect 314782 384618 314866 384854
rect 315102 384618 334546 384854
rect 334782 384618 334866 384854
rect 335102 384618 354546 384854
rect 354782 384618 354866 384854
rect 355102 384618 374546 384854
rect 374782 384618 374866 384854
rect 375102 384618 394546 384854
rect 394782 384618 394866 384854
rect 395102 384618 414546 384854
rect 414782 384618 414866 384854
rect 415102 384618 434546 384854
rect 434782 384618 434866 384854
rect 435102 384618 454546 384854
rect 454782 384618 454866 384854
rect 455102 384618 474546 384854
rect 474782 384618 474866 384854
rect 475102 384618 494546 384854
rect 494782 384618 494866 384854
rect 495102 384618 514546 384854
rect 514782 384618 514866 384854
rect 515102 384618 534546 384854
rect 534782 384618 534866 384854
rect 535102 384618 554546 384854
rect 554782 384618 554866 384854
rect 555102 384618 574546 384854
rect 574782 384618 574866 384854
rect 575102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 10826 381454
rect 11062 381218 11146 381454
rect 11382 381218 30826 381454
rect 31062 381218 31146 381454
rect 31382 381218 50826 381454
rect 51062 381218 51146 381454
rect 51382 381218 70826 381454
rect 71062 381218 71146 381454
rect 71382 381218 90826 381454
rect 91062 381218 91146 381454
rect 91382 381218 110826 381454
rect 111062 381218 111146 381454
rect 111382 381218 130826 381454
rect 131062 381218 131146 381454
rect 131382 381218 150826 381454
rect 151062 381218 151146 381454
rect 151382 381218 170826 381454
rect 171062 381218 171146 381454
rect 171382 381218 190826 381454
rect 191062 381218 191146 381454
rect 191382 381218 210826 381454
rect 211062 381218 211146 381454
rect 211382 381218 230826 381454
rect 231062 381218 231146 381454
rect 231382 381218 250826 381454
rect 251062 381218 251146 381454
rect 251382 381218 270826 381454
rect 271062 381218 271146 381454
rect 271382 381218 290826 381454
rect 291062 381218 291146 381454
rect 291382 381218 310826 381454
rect 311062 381218 311146 381454
rect 311382 381218 330826 381454
rect 331062 381218 331146 381454
rect 331382 381218 350826 381454
rect 351062 381218 351146 381454
rect 351382 381218 370826 381454
rect 371062 381218 371146 381454
rect 371382 381218 390826 381454
rect 391062 381218 391146 381454
rect 391382 381218 410826 381454
rect 411062 381218 411146 381454
rect 411382 381218 430826 381454
rect 431062 381218 431146 381454
rect 431382 381218 450826 381454
rect 451062 381218 451146 381454
rect 451382 381218 470826 381454
rect 471062 381218 471146 381454
rect 471382 381218 490826 381454
rect 491062 381218 491146 381454
rect 491382 381218 510826 381454
rect 511062 381218 511146 381454
rect 511382 381218 530826 381454
rect 531062 381218 531146 381454
rect 531382 381218 550826 381454
rect 551062 381218 551146 381454
rect 551382 381218 570826 381454
rect 571062 381218 571146 381454
rect 571382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 10826 381134
rect 11062 380898 11146 381134
rect 11382 380898 30826 381134
rect 31062 380898 31146 381134
rect 31382 380898 50826 381134
rect 51062 380898 51146 381134
rect 51382 380898 70826 381134
rect 71062 380898 71146 381134
rect 71382 380898 90826 381134
rect 91062 380898 91146 381134
rect 91382 380898 110826 381134
rect 111062 380898 111146 381134
rect 111382 380898 130826 381134
rect 131062 380898 131146 381134
rect 131382 380898 150826 381134
rect 151062 380898 151146 381134
rect 151382 380898 170826 381134
rect 171062 380898 171146 381134
rect 171382 380898 190826 381134
rect 191062 380898 191146 381134
rect 191382 380898 210826 381134
rect 211062 380898 211146 381134
rect 211382 380898 230826 381134
rect 231062 380898 231146 381134
rect 231382 380898 250826 381134
rect 251062 380898 251146 381134
rect 251382 380898 270826 381134
rect 271062 380898 271146 381134
rect 271382 380898 290826 381134
rect 291062 380898 291146 381134
rect 291382 380898 310826 381134
rect 311062 380898 311146 381134
rect 311382 380898 330826 381134
rect 331062 380898 331146 381134
rect 331382 380898 350826 381134
rect 351062 380898 351146 381134
rect 351382 380898 370826 381134
rect 371062 380898 371146 381134
rect 371382 380898 390826 381134
rect 391062 380898 391146 381134
rect 391382 380898 410826 381134
rect 411062 380898 411146 381134
rect 411382 380898 430826 381134
rect 431062 380898 431146 381134
rect 431382 380898 450826 381134
rect 451062 380898 451146 381134
rect 451382 380898 470826 381134
rect 471062 380898 471146 381134
rect 471382 380898 490826 381134
rect 491062 380898 491146 381134
rect 491382 380898 510826 381134
rect 511062 380898 511146 381134
rect 511382 380898 530826 381134
rect 531062 380898 531146 381134
rect 531382 380898 550826 381134
rect 551062 380898 551146 381134
rect 551382 380898 570826 381134
rect 571062 380898 571146 381134
rect 571382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 11986 374614
rect 12222 374378 12306 374614
rect 12542 374378 31986 374614
rect 32222 374378 32306 374614
rect 32542 374378 51986 374614
rect 52222 374378 52306 374614
rect 52542 374378 71986 374614
rect 72222 374378 72306 374614
rect 72542 374378 91986 374614
rect 92222 374378 92306 374614
rect 92542 374378 111986 374614
rect 112222 374378 112306 374614
rect 112542 374378 131986 374614
rect 132222 374378 132306 374614
rect 132542 374378 151986 374614
rect 152222 374378 152306 374614
rect 152542 374378 171986 374614
rect 172222 374378 172306 374614
rect 172542 374378 191986 374614
rect 192222 374378 192306 374614
rect 192542 374378 211986 374614
rect 212222 374378 212306 374614
rect 212542 374378 231986 374614
rect 232222 374378 232306 374614
rect 232542 374378 251986 374614
rect 252222 374378 252306 374614
rect 252542 374378 271986 374614
rect 272222 374378 272306 374614
rect 272542 374378 291986 374614
rect 292222 374378 292306 374614
rect 292542 374378 311986 374614
rect 312222 374378 312306 374614
rect 312542 374378 331986 374614
rect 332222 374378 332306 374614
rect 332542 374378 351986 374614
rect 352222 374378 352306 374614
rect 352542 374378 371986 374614
rect 372222 374378 372306 374614
rect 372542 374378 391986 374614
rect 392222 374378 392306 374614
rect 392542 374378 411986 374614
rect 412222 374378 412306 374614
rect 412542 374378 431986 374614
rect 432222 374378 432306 374614
rect 432542 374378 451986 374614
rect 452222 374378 452306 374614
rect 452542 374378 471986 374614
rect 472222 374378 472306 374614
rect 472542 374378 491986 374614
rect 492222 374378 492306 374614
rect 492542 374378 511986 374614
rect 512222 374378 512306 374614
rect 512542 374378 531986 374614
rect 532222 374378 532306 374614
rect 532542 374378 551986 374614
rect 552222 374378 552306 374614
rect 552542 374378 571986 374614
rect 572222 374378 572306 374614
rect 572542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 11986 374294
rect 12222 374058 12306 374294
rect 12542 374058 31986 374294
rect 32222 374058 32306 374294
rect 32542 374058 51986 374294
rect 52222 374058 52306 374294
rect 52542 374058 71986 374294
rect 72222 374058 72306 374294
rect 72542 374058 91986 374294
rect 92222 374058 92306 374294
rect 92542 374058 111986 374294
rect 112222 374058 112306 374294
rect 112542 374058 131986 374294
rect 132222 374058 132306 374294
rect 132542 374058 151986 374294
rect 152222 374058 152306 374294
rect 152542 374058 171986 374294
rect 172222 374058 172306 374294
rect 172542 374058 191986 374294
rect 192222 374058 192306 374294
rect 192542 374058 211986 374294
rect 212222 374058 212306 374294
rect 212542 374058 231986 374294
rect 232222 374058 232306 374294
rect 232542 374058 251986 374294
rect 252222 374058 252306 374294
rect 252542 374058 271986 374294
rect 272222 374058 272306 374294
rect 272542 374058 291986 374294
rect 292222 374058 292306 374294
rect 292542 374058 311986 374294
rect 312222 374058 312306 374294
rect 312542 374058 331986 374294
rect 332222 374058 332306 374294
rect 332542 374058 351986 374294
rect 352222 374058 352306 374294
rect 352542 374058 371986 374294
rect 372222 374058 372306 374294
rect 372542 374058 391986 374294
rect 392222 374058 392306 374294
rect 392542 374058 411986 374294
rect 412222 374058 412306 374294
rect 412542 374058 431986 374294
rect 432222 374058 432306 374294
rect 432542 374058 451986 374294
rect 452222 374058 452306 374294
rect 452542 374058 471986 374294
rect 472222 374058 472306 374294
rect 472542 374058 491986 374294
rect 492222 374058 492306 374294
rect 492542 374058 511986 374294
rect 512222 374058 512306 374294
rect 512542 374058 531986 374294
rect 532222 374058 532306 374294
rect 532542 374058 551986 374294
rect 552222 374058 552306 374294
rect 552542 374058 571986 374294
rect 572222 374058 572306 374294
rect 572542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 8266 370894
rect 8502 370658 8586 370894
rect 8822 370658 28266 370894
rect 28502 370658 28586 370894
rect 28822 370658 48266 370894
rect 48502 370658 48586 370894
rect 48822 370658 68266 370894
rect 68502 370658 68586 370894
rect 68822 370658 88266 370894
rect 88502 370658 88586 370894
rect 88822 370658 108266 370894
rect 108502 370658 108586 370894
rect 108822 370658 128266 370894
rect 128502 370658 128586 370894
rect 128822 370658 148266 370894
rect 148502 370658 148586 370894
rect 148822 370658 168266 370894
rect 168502 370658 168586 370894
rect 168822 370658 188266 370894
rect 188502 370658 188586 370894
rect 188822 370658 208266 370894
rect 208502 370658 208586 370894
rect 208822 370658 228266 370894
rect 228502 370658 228586 370894
rect 228822 370658 248266 370894
rect 248502 370658 248586 370894
rect 248822 370658 268266 370894
rect 268502 370658 268586 370894
rect 268822 370658 288266 370894
rect 288502 370658 288586 370894
rect 288822 370658 308266 370894
rect 308502 370658 308586 370894
rect 308822 370658 328266 370894
rect 328502 370658 328586 370894
rect 328822 370658 348266 370894
rect 348502 370658 348586 370894
rect 348822 370658 368266 370894
rect 368502 370658 368586 370894
rect 368822 370658 388266 370894
rect 388502 370658 388586 370894
rect 388822 370658 408266 370894
rect 408502 370658 408586 370894
rect 408822 370658 428266 370894
rect 428502 370658 428586 370894
rect 428822 370658 448266 370894
rect 448502 370658 448586 370894
rect 448822 370658 468266 370894
rect 468502 370658 468586 370894
rect 468822 370658 488266 370894
rect 488502 370658 488586 370894
rect 488822 370658 508266 370894
rect 508502 370658 508586 370894
rect 508822 370658 528266 370894
rect 528502 370658 528586 370894
rect 528822 370658 548266 370894
rect 548502 370658 548586 370894
rect 548822 370658 568266 370894
rect 568502 370658 568586 370894
rect 568822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 8266 370574
rect 8502 370338 8586 370574
rect 8822 370338 28266 370574
rect 28502 370338 28586 370574
rect 28822 370338 48266 370574
rect 48502 370338 48586 370574
rect 48822 370338 68266 370574
rect 68502 370338 68586 370574
rect 68822 370338 88266 370574
rect 88502 370338 88586 370574
rect 88822 370338 108266 370574
rect 108502 370338 108586 370574
rect 108822 370338 128266 370574
rect 128502 370338 128586 370574
rect 128822 370338 148266 370574
rect 148502 370338 148586 370574
rect 148822 370338 168266 370574
rect 168502 370338 168586 370574
rect 168822 370338 188266 370574
rect 188502 370338 188586 370574
rect 188822 370338 208266 370574
rect 208502 370338 208586 370574
rect 208822 370338 228266 370574
rect 228502 370338 228586 370574
rect 228822 370338 248266 370574
rect 248502 370338 248586 370574
rect 248822 370338 268266 370574
rect 268502 370338 268586 370574
rect 268822 370338 288266 370574
rect 288502 370338 288586 370574
rect 288822 370338 308266 370574
rect 308502 370338 308586 370574
rect 308822 370338 328266 370574
rect 328502 370338 328586 370574
rect 328822 370338 348266 370574
rect 348502 370338 348586 370574
rect 348822 370338 368266 370574
rect 368502 370338 368586 370574
rect 368822 370338 388266 370574
rect 388502 370338 388586 370574
rect 388822 370338 408266 370574
rect 408502 370338 408586 370574
rect 408822 370338 428266 370574
rect 428502 370338 428586 370574
rect 428822 370338 448266 370574
rect 448502 370338 448586 370574
rect 448822 370338 468266 370574
rect 468502 370338 468586 370574
rect 468822 370338 488266 370574
rect 488502 370338 488586 370574
rect 488822 370338 508266 370574
rect 508502 370338 508586 370574
rect 508822 370338 528266 370574
rect 528502 370338 528586 370574
rect 528822 370338 548266 370574
rect 548502 370338 548586 370574
rect 548822 370338 568266 370574
rect 568502 370338 568586 370574
rect 568822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 4546 367174
rect 4782 366938 4866 367174
rect 5102 366938 24546 367174
rect 24782 366938 24866 367174
rect 25102 366938 44546 367174
rect 44782 366938 44866 367174
rect 45102 366938 64546 367174
rect 64782 366938 64866 367174
rect 65102 366938 84546 367174
rect 84782 366938 84866 367174
rect 85102 366938 104546 367174
rect 104782 366938 104866 367174
rect 105102 366938 124546 367174
rect 124782 366938 124866 367174
rect 125102 366938 144546 367174
rect 144782 366938 144866 367174
rect 145102 366938 164546 367174
rect 164782 366938 164866 367174
rect 165102 366938 184546 367174
rect 184782 366938 184866 367174
rect 185102 366938 204546 367174
rect 204782 366938 204866 367174
rect 205102 366938 224546 367174
rect 224782 366938 224866 367174
rect 225102 366938 244546 367174
rect 244782 366938 244866 367174
rect 245102 366938 264546 367174
rect 264782 366938 264866 367174
rect 265102 366938 284546 367174
rect 284782 366938 284866 367174
rect 285102 366938 304546 367174
rect 304782 366938 304866 367174
rect 305102 366938 324546 367174
rect 324782 366938 324866 367174
rect 325102 366938 344546 367174
rect 344782 366938 344866 367174
rect 345102 366938 364546 367174
rect 364782 366938 364866 367174
rect 365102 366938 384546 367174
rect 384782 366938 384866 367174
rect 385102 366938 404546 367174
rect 404782 366938 404866 367174
rect 405102 366938 424546 367174
rect 424782 366938 424866 367174
rect 425102 366938 444546 367174
rect 444782 366938 444866 367174
rect 445102 366938 464546 367174
rect 464782 366938 464866 367174
rect 465102 366938 484546 367174
rect 484782 366938 484866 367174
rect 485102 366938 504546 367174
rect 504782 366938 504866 367174
rect 505102 366938 524546 367174
rect 524782 366938 524866 367174
rect 525102 366938 544546 367174
rect 544782 366938 544866 367174
rect 545102 366938 564546 367174
rect 564782 366938 564866 367174
rect 565102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 4546 366854
rect 4782 366618 4866 366854
rect 5102 366618 24546 366854
rect 24782 366618 24866 366854
rect 25102 366618 44546 366854
rect 44782 366618 44866 366854
rect 45102 366618 64546 366854
rect 64782 366618 64866 366854
rect 65102 366618 84546 366854
rect 84782 366618 84866 366854
rect 85102 366618 104546 366854
rect 104782 366618 104866 366854
rect 105102 366618 124546 366854
rect 124782 366618 124866 366854
rect 125102 366618 144546 366854
rect 144782 366618 144866 366854
rect 145102 366618 164546 366854
rect 164782 366618 164866 366854
rect 165102 366618 184546 366854
rect 184782 366618 184866 366854
rect 185102 366618 204546 366854
rect 204782 366618 204866 366854
rect 205102 366618 224546 366854
rect 224782 366618 224866 366854
rect 225102 366618 244546 366854
rect 244782 366618 244866 366854
rect 245102 366618 264546 366854
rect 264782 366618 264866 366854
rect 265102 366618 284546 366854
rect 284782 366618 284866 366854
rect 285102 366618 304546 366854
rect 304782 366618 304866 366854
rect 305102 366618 324546 366854
rect 324782 366618 324866 366854
rect 325102 366618 344546 366854
rect 344782 366618 344866 366854
rect 345102 366618 364546 366854
rect 364782 366618 364866 366854
rect 365102 366618 384546 366854
rect 384782 366618 384866 366854
rect 385102 366618 404546 366854
rect 404782 366618 404866 366854
rect 405102 366618 424546 366854
rect 424782 366618 424866 366854
rect 425102 366618 444546 366854
rect 444782 366618 444866 366854
rect 445102 366618 464546 366854
rect 464782 366618 464866 366854
rect 465102 366618 484546 366854
rect 484782 366618 484866 366854
rect 485102 366618 504546 366854
rect 504782 366618 504866 366854
rect 505102 366618 524546 366854
rect 524782 366618 524866 366854
rect 525102 366618 544546 366854
rect 544782 366618 544866 366854
rect 545102 366618 564546 366854
rect 564782 366618 564866 366854
rect 565102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 826 363454
rect 1062 363218 1146 363454
rect 1382 363218 20826 363454
rect 21062 363218 21146 363454
rect 21382 363218 40826 363454
rect 41062 363218 41146 363454
rect 41382 363218 60826 363454
rect 61062 363218 61146 363454
rect 61382 363218 80826 363454
rect 81062 363218 81146 363454
rect 81382 363218 100826 363454
rect 101062 363218 101146 363454
rect 101382 363218 120826 363454
rect 121062 363218 121146 363454
rect 121382 363218 140826 363454
rect 141062 363218 141146 363454
rect 141382 363218 160826 363454
rect 161062 363218 161146 363454
rect 161382 363218 180826 363454
rect 181062 363218 181146 363454
rect 181382 363218 200826 363454
rect 201062 363218 201146 363454
rect 201382 363218 220826 363454
rect 221062 363218 221146 363454
rect 221382 363218 240826 363454
rect 241062 363218 241146 363454
rect 241382 363218 260826 363454
rect 261062 363218 261146 363454
rect 261382 363218 280826 363454
rect 281062 363218 281146 363454
rect 281382 363218 300826 363454
rect 301062 363218 301146 363454
rect 301382 363218 320826 363454
rect 321062 363218 321146 363454
rect 321382 363218 340826 363454
rect 341062 363218 341146 363454
rect 341382 363218 360826 363454
rect 361062 363218 361146 363454
rect 361382 363218 380826 363454
rect 381062 363218 381146 363454
rect 381382 363218 400826 363454
rect 401062 363218 401146 363454
rect 401382 363218 420826 363454
rect 421062 363218 421146 363454
rect 421382 363218 440826 363454
rect 441062 363218 441146 363454
rect 441382 363218 460826 363454
rect 461062 363218 461146 363454
rect 461382 363218 480826 363454
rect 481062 363218 481146 363454
rect 481382 363218 500826 363454
rect 501062 363218 501146 363454
rect 501382 363218 520826 363454
rect 521062 363218 521146 363454
rect 521382 363218 540826 363454
rect 541062 363218 541146 363454
rect 541382 363218 560826 363454
rect 561062 363218 561146 363454
rect 561382 363218 580826 363454
rect 581062 363218 581146 363454
rect 581382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 826 363134
rect 1062 362898 1146 363134
rect 1382 362898 20826 363134
rect 21062 362898 21146 363134
rect 21382 362898 40826 363134
rect 41062 362898 41146 363134
rect 41382 362898 60826 363134
rect 61062 362898 61146 363134
rect 61382 362898 80826 363134
rect 81062 362898 81146 363134
rect 81382 362898 100826 363134
rect 101062 362898 101146 363134
rect 101382 362898 120826 363134
rect 121062 362898 121146 363134
rect 121382 362898 140826 363134
rect 141062 362898 141146 363134
rect 141382 362898 160826 363134
rect 161062 362898 161146 363134
rect 161382 362898 180826 363134
rect 181062 362898 181146 363134
rect 181382 362898 200826 363134
rect 201062 362898 201146 363134
rect 201382 362898 220826 363134
rect 221062 362898 221146 363134
rect 221382 362898 240826 363134
rect 241062 362898 241146 363134
rect 241382 362898 260826 363134
rect 261062 362898 261146 363134
rect 261382 362898 280826 363134
rect 281062 362898 281146 363134
rect 281382 362898 300826 363134
rect 301062 362898 301146 363134
rect 301382 362898 320826 363134
rect 321062 362898 321146 363134
rect 321382 362898 340826 363134
rect 341062 362898 341146 363134
rect 341382 362898 360826 363134
rect 361062 362898 361146 363134
rect 361382 362898 380826 363134
rect 381062 362898 381146 363134
rect 381382 362898 400826 363134
rect 401062 362898 401146 363134
rect 401382 362898 420826 363134
rect 421062 362898 421146 363134
rect 421382 362898 440826 363134
rect 441062 362898 441146 363134
rect 441382 362898 460826 363134
rect 461062 362898 461146 363134
rect 461382 362898 480826 363134
rect 481062 362898 481146 363134
rect 481382 362898 500826 363134
rect 501062 362898 501146 363134
rect 501382 362898 520826 363134
rect 521062 362898 521146 363134
rect 521382 362898 540826 363134
rect 541062 362898 541146 363134
rect 541382 362898 560826 363134
rect 561062 362898 561146 363134
rect 561382 362898 580826 363134
rect 581062 362898 581146 363134
rect 581382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 21986 356614
rect 22222 356378 22306 356614
rect 22542 356378 41986 356614
rect 42222 356378 42306 356614
rect 42542 356378 61986 356614
rect 62222 356378 62306 356614
rect 62542 356378 81986 356614
rect 82222 356378 82306 356614
rect 82542 356378 101986 356614
rect 102222 356378 102306 356614
rect 102542 356378 121986 356614
rect 122222 356378 122306 356614
rect 122542 356378 141986 356614
rect 142222 356378 142306 356614
rect 142542 356378 161986 356614
rect 162222 356378 162306 356614
rect 162542 356378 181986 356614
rect 182222 356378 182306 356614
rect 182542 356378 201986 356614
rect 202222 356378 202306 356614
rect 202542 356378 221986 356614
rect 222222 356378 222306 356614
rect 222542 356378 241986 356614
rect 242222 356378 242306 356614
rect 242542 356378 261986 356614
rect 262222 356378 262306 356614
rect 262542 356378 281986 356614
rect 282222 356378 282306 356614
rect 282542 356378 301986 356614
rect 302222 356378 302306 356614
rect 302542 356378 321986 356614
rect 322222 356378 322306 356614
rect 322542 356378 341986 356614
rect 342222 356378 342306 356614
rect 342542 356378 361986 356614
rect 362222 356378 362306 356614
rect 362542 356378 381986 356614
rect 382222 356378 382306 356614
rect 382542 356378 401986 356614
rect 402222 356378 402306 356614
rect 402542 356378 421986 356614
rect 422222 356378 422306 356614
rect 422542 356378 441986 356614
rect 442222 356378 442306 356614
rect 442542 356378 461986 356614
rect 462222 356378 462306 356614
rect 462542 356378 481986 356614
rect 482222 356378 482306 356614
rect 482542 356378 501986 356614
rect 502222 356378 502306 356614
rect 502542 356378 521986 356614
rect 522222 356378 522306 356614
rect 522542 356378 541986 356614
rect 542222 356378 542306 356614
rect 542542 356378 561986 356614
rect 562222 356378 562306 356614
rect 562542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 21986 356294
rect 22222 356058 22306 356294
rect 22542 356058 41986 356294
rect 42222 356058 42306 356294
rect 42542 356058 61986 356294
rect 62222 356058 62306 356294
rect 62542 356058 81986 356294
rect 82222 356058 82306 356294
rect 82542 356058 101986 356294
rect 102222 356058 102306 356294
rect 102542 356058 121986 356294
rect 122222 356058 122306 356294
rect 122542 356058 141986 356294
rect 142222 356058 142306 356294
rect 142542 356058 161986 356294
rect 162222 356058 162306 356294
rect 162542 356058 181986 356294
rect 182222 356058 182306 356294
rect 182542 356058 201986 356294
rect 202222 356058 202306 356294
rect 202542 356058 221986 356294
rect 222222 356058 222306 356294
rect 222542 356058 241986 356294
rect 242222 356058 242306 356294
rect 242542 356058 261986 356294
rect 262222 356058 262306 356294
rect 262542 356058 281986 356294
rect 282222 356058 282306 356294
rect 282542 356058 301986 356294
rect 302222 356058 302306 356294
rect 302542 356058 321986 356294
rect 322222 356058 322306 356294
rect 322542 356058 341986 356294
rect 342222 356058 342306 356294
rect 342542 356058 361986 356294
rect 362222 356058 362306 356294
rect 362542 356058 381986 356294
rect 382222 356058 382306 356294
rect 382542 356058 401986 356294
rect 402222 356058 402306 356294
rect 402542 356058 421986 356294
rect 422222 356058 422306 356294
rect 422542 356058 441986 356294
rect 442222 356058 442306 356294
rect 442542 356058 461986 356294
rect 462222 356058 462306 356294
rect 462542 356058 481986 356294
rect 482222 356058 482306 356294
rect 482542 356058 501986 356294
rect 502222 356058 502306 356294
rect 502542 356058 521986 356294
rect 522222 356058 522306 356294
rect 522542 356058 541986 356294
rect 542222 356058 542306 356294
rect 542542 356058 561986 356294
rect 562222 356058 562306 356294
rect 562542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 18266 352894
rect 18502 352658 18586 352894
rect 18822 352658 38266 352894
rect 38502 352658 38586 352894
rect 38822 352658 58266 352894
rect 58502 352658 58586 352894
rect 58822 352658 78266 352894
rect 78502 352658 78586 352894
rect 78822 352658 98266 352894
rect 98502 352658 98586 352894
rect 98822 352658 118266 352894
rect 118502 352658 118586 352894
rect 118822 352658 138266 352894
rect 138502 352658 138586 352894
rect 138822 352658 158266 352894
rect 158502 352658 158586 352894
rect 158822 352658 178266 352894
rect 178502 352658 178586 352894
rect 178822 352658 198266 352894
rect 198502 352658 198586 352894
rect 198822 352658 218266 352894
rect 218502 352658 218586 352894
rect 218822 352658 238266 352894
rect 238502 352658 238586 352894
rect 238822 352658 258266 352894
rect 258502 352658 258586 352894
rect 258822 352658 278266 352894
rect 278502 352658 278586 352894
rect 278822 352658 298266 352894
rect 298502 352658 298586 352894
rect 298822 352658 318266 352894
rect 318502 352658 318586 352894
rect 318822 352658 338266 352894
rect 338502 352658 338586 352894
rect 338822 352658 358266 352894
rect 358502 352658 358586 352894
rect 358822 352658 378266 352894
rect 378502 352658 378586 352894
rect 378822 352658 398266 352894
rect 398502 352658 398586 352894
rect 398822 352658 418266 352894
rect 418502 352658 418586 352894
rect 418822 352658 438266 352894
rect 438502 352658 438586 352894
rect 438822 352658 458266 352894
rect 458502 352658 458586 352894
rect 458822 352658 478266 352894
rect 478502 352658 478586 352894
rect 478822 352658 498266 352894
rect 498502 352658 498586 352894
rect 498822 352658 518266 352894
rect 518502 352658 518586 352894
rect 518822 352658 538266 352894
rect 538502 352658 538586 352894
rect 538822 352658 558266 352894
rect 558502 352658 558586 352894
rect 558822 352658 578266 352894
rect 578502 352658 578586 352894
rect 578822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 18266 352574
rect 18502 352338 18586 352574
rect 18822 352338 38266 352574
rect 38502 352338 38586 352574
rect 38822 352338 58266 352574
rect 58502 352338 58586 352574
rect 58822 352338 78266 352574
rect 78502 352338 78586 352574
rect 78822 352338 98266 352574
rect 98502 352338 98586 352574
rect 98822 352338 118266 352574
rect 118502 352338 118586 352574
rect 118822 352338 138266 352574
rect 138502 352338 138586 352574
rect 138822 352338 158266 352574
rect 158502 352338 158586 352574
rect 158822 352338 178266 352574
rect 178502 352338 178586 352574
rect 178822 352338 198266 352574
rect 198502 352338 198586 352574
rect 198822 352338 218266 352574
rect 218502 352338 218586 352574
rect 218822 352338 238266 352574
rect 238502 352338 238586 352574
rect 238822 352338 258266 352574
rect 258502 352338 258586 352574
rect 258822 352338 278266 352574
rect 278502 352338 278586 352574
rect 278822 352338 298266 352574
rect 298502 352338 298586 352574
rect 298822 352338 318266 352574
rect 318502 352338 318586 352574
rect 318822 352338 338266 352574
rect 338502 352338 338586 352574
rect 338822 352338 358266 352574
rect 358502 352338 358586 352574
rect 358822 352338 378266 352574
rect 378502 352338 378586 352574
rect 378822 352338 398266 352574
rect 398502 352338 398586 352574
rect 398822 352338 418266 352574
rect 418502 352338 418586 352574
rect 418822 352338 438266 352574
rect 438502 352338 438586 352574
rect 438822 352338 458266 352574
rect 458502 352338 458586 352574
rect 458822 352338 478266 352574
rect 478502 352338 478586 352574
rect 478822 352338 498266 352574
rect 498502 352338 498586 352574
rect 498822 352338 518266 352574
rect 518502 352338 518586 352574
rect 518822 352338 538266 352574
rect 538502 352338 538586 352574
rect 538822 352338 558266 352574
rect 558502 352338 558586 352574
rect 558822 352338 578266 352574
rect 578502 352338 578586 352574
rect 578822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 14546 349174
rect 14782 348938 14866 349174
rect 15102 348938 34546 349174
rect 34782 348938 34866 349174
rect 35102 348938 54546 349174
rect 54782 348938 54866 349174
rect 55102 348938 74546 349174
rect 74782 348938 74866 349174
rect 75102 348938 94546 349174
rect 94782 348938 94866 349174
rect 95102 348938 114546 349174
rect 114782 348938 114866 349174
rect 115102 348938 134546 349174
rect 134782 348938 134866 349174
rect 135102 348938 154546 349174
rect 154782 348938 154866 349174
rect 155102 348938 174546 349174
rect 174782 348938 174866 349174
rect 175102 348938 194546 349174
rect 194782 348938 194866 349174
rect 195102 348938 214546 349174
rect 214782 348938 214866 349174
rect 215102 348938 234546 349174
rect 234782 348938 234866 349174
rect 235102 348938 254546 349174
rect 254782 348938 254866 349174
rect 255102 348938 274546 349174
rect 274782 348938 274866 349174
rect 275102 348938 294546 349174
rect 294782 348938 294866 349174
rect 295102 348938 314546 349174
rect 314782 348938 314866 349174
rect 315102 348938 334546 349174
rect 334782 348938 334866 349174
rect 335102 348938 354546 349174
rect 354782 348938 354866 349174
rect 355102 348938 374546 349174
rect 374782 348938 374866 349174
rect 375102 348938 394546 349174
rect 394782 348938 394866 349174
rect 395102 348938 414546 349174
rect 414782 348938 414866 349174
rect 415102 348938 434546 349174
rect 434782 348938 434866 349174
rect 435102 348938 454546 349174
rect 454782 348938 454866 349174
rect 455102 348938 474546 349174
rect 474782 348938 474866 349174
rect 475102 348938 494546 349174
rect 494782 348938 494866 349174
rect 495102 348938 514546 349174
rect 514782 348938 514866 349174
rect 515102 348938 534546 349174
rect 534782 348938 534866 349174
rect 535102 348938 554546 349174
rect 554782 348938 554866 349174
rect 555102 348938 574546 349174
rect 574782 348938 574866 349174
rect 575102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 14546 348854
rect 14782 348618 14866 348854
rect 15102 348618 34546 348854
rect 34782 348618 34866 348854
rect 35102 348618 54546 348854
rect 54782 348618 54866 348854
rect 55102 348618 74546 348854
rect 74782 348618 74866 348854
rect 75102 348618 94546 348854
rect 94782 348618 94866 348854
rect 95102 348618 114546 348854
rect 114782 348618 114866 348854
rect 115102 348618 134546 348854
rect 134782 348618 134866 348854
rect 135102 348618 154546 348854
rect 154782 348618 154866 348854
rect 155102 348618 174546 348854
rect 174782 348618 174866 348854
rect 175102 348618 194546 348854
rect 194782 348618 194866 348854
rect 195102 348618 214546 348854
rect 214782 348618 214866 348854
rect 215102 348618 234546 348854
rect 234782 348618 234866 348854
rect 235102 348618 254546 348854
rect 254782 348618 254866 348854
rect 255102 348618 274546 348854
rect 274782 348618 274866 348854
rect 275102 348618 294546 348854
rect 294782 348618 294866 348854
rect 295102 348618 314546 348854
rect 314782 348618 314866 348854
rect 315102 348618 334546 348854
rect 334782 348618 334866 348854
rect 335102 348618 354546 348854
rect 354782 348618 354866 348854
rect 355102 348618 374546 348854
rect 374782 348618 374866 348854
rect 375102 348618 394546 348854
rect 394782 348618 394866 348854
rect 395102 348618 414546 348854
rect 414782 348618 414866 348854
rect 415102 348618 434546 348854
rect 434782 348618 434866 348854
rect 435102 348618 454546 348854
rect 454782 348618 454866 348854
rect 455102 348618 474546 348854
rect 474782 348618 474866 348854
rect 475102 348618 494546 348854
rect 494782 348618 494866 348854
rect 495102 348618 514546 348854
rect 514782 348618 514866 348854
rect 515102 348618 534546 348854
rect 534782 348618 534866 348854
rect 535102 348618 554546 348854
rect 554782 348618 554866 348854
rect 555102 348618 574546 348854
rect 574782 348618 574866 348854
rect 575102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 10826 345454
rect 11062 345218 11146 345454
rect 11382 345218 30826 345454
rect 31062 345218 31146 345454
rect 31382 345218 50826 345454
rect 51062 345218 51146 345454
rect 51382 345218 70826 345454
rect 71062 345218 71146 345454
rect 71382 345218 90826 345454
rect 91062 345218 91146 345454
rect 91382 345218 110826 345454
rect 111062 345218 111146 345454
rect 111382 345218 130826 345454
rect 131062 345218 131146 345454
rect 131382 345218 150826 345454
rect 151062 345218 151146 345454
rect 151382 345218 170826 345454
rect 171062 345218 171146 345454
rect 171382 345218 190826 345454
rect 191062 345218 191146 345454
rect 191382 345218 210826 345454
rect 211062 345218 211146 345454
rect 211382 345218 230826 345454
rect 231062 345218 231146 345454
rect 231382 345218 250826 345454
rect 251062 345218 251146 345454
rect 251382 345218 270826 345454
rect 271062 345218 271146 345454
rect 271382 345218 290826 345454
rect 291062 345218 291146 345454
rect 291382 345218 310826 345454
rect 311062 345218 311146 345454
rect 311382 345218 330826 345454
rect 331062 345218 331146 345454
rect 331382 345218 350826 345454
rect 351062 345218 351146 345454
rect 351382 345218 370826 345454
rect 371062 345218 371146 345454
rect 371382 345218 390826 345454
rect 391062 345218 391146 345454
rect 391382 345218 410826 345454
rect 411062 345218 411146 345454
rect 411382 345218 430826 345454
rect 431062 345218 431146 345454
rect 431382 345218 450826 345454
rect 451062 345218 451146 345454
rect 451382 345218 470826 345454
rect 471062 345218 471146 345454
rect 471382 345218 490826 345454
rect 491062 345218 491146 345454
rect 491382 345218 510826 345454
rect 511062 345218 511146 345454
rect 511382 345218 530826 345454
rect 531062 345218 531146 345454
rect 531382 345218 550826 345454
rect 551062 345218 551146 345454
rect 551382 345218 570826 345454
rect 571062 345218 571146 345454
rect 571382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 10826 345134
rect 11062 344898 11146 345134
rect 11382 344898 30826 345134
rect 31062 344898 31146 345134
rect 31382 344898 50826 345134
rect 51062 344898 51146 345134
rect 51382 344898 70826 345134
rect 71062 344898 71146 345134
rect 71382 344898 90826 345134
rect 91062 344898 91146 345134
rect 91382 344898 110826 345134
rect 111062 344898 111146 345134
rect 111382 344898 130826 345134
rect 131062 344898 131146 345134
rect 131382 344898 150826 345134
rect 151062 344898 151146 345134
rect 151382 344898 170826 345134
rect 171062 344898 171146 345134
rect 171382 344898 190826 345134
rect 191062 344898 191146 345134
rect 191382 344898 210826 345134
rect 211062 344898 211146 345134
rect 211382 344898 230826 345134
rect 231062 344898 231146 345134
rect 231382 344898 250826 345134
rect 251062 344898 251146 345134
rect 251382 344898 270826 345134
rect 271062 344898 271146 345134
rect 271382 344898 290826 345134
rect 291062 344898 291146 345134
rect 291382 344898 310826 345134
rect 311062 344898 311146 345134
rect 311382 344898 330826 345134
rect 331062 344898 331146 345134
rect 331382 344898 350826 345134
rect 351062 344898 351146 345134
rect 351382 344898 370826 345134
rect 371062 344898 371146 345134
rect 371382 344898 390826 345134
rect 391062 344898 391146 345134
rect 391382 344898 410826 345134
rect 411062 344898 411146 345134
rect 411382 344898 430826 345134
rect 431062 344898 431146 345134
rect 431382 344898 450826 345134
rect 451062 344898 451146 345134
rect 451382 344898 470826 345134
rect 471062 344898 471146 345134
rect 471382 344898 490826 345134
rect 491062 344898 491146 345134
rect 491382 344898 510826 345134
rect 511062 344898 511146 345134
rect 511382 344898 530826 345134
rect 531062 344898 531146 345134
rect 531382 344898 550826 345134
rect 551062 344898 551146 345134
rect 551382 344898 570826 345134
rect 571062 344898 571146 345134
rect 571382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 11986 338614
rect 12222 338378 12306 338614
rect 12542 338378 31986 338614
rect 32222 338378 32306 338614
rect 32542 338378 51986 338614
rect 52222 338378 52306 338614
rect 52542 338378 71986 338614
rect 72222 338378 72306 338614
rect 72542 338378 91986 338614
rect 92222 338378 92306 338614
rect 92542 338378 111986 338614
rect 112222 338378 112306 338614
rect 112542 338378 131986 338614
rect 132222 338378 132306 338614
rect 132542 338378 151986 338614
rect 152222 338378 152306 338614
rect 152542 338378 171986 338614
rect 172222 338378 172306 338614
rect 172542 338378 191986 338614
rect 192222 338378 192306 338614
rect 192542 338378 211986 338614
rect 212222 338378 212306 338614
rect 212542 338378 231986 338614
rect 232222 338378 232306 338614
rect 232542 338378 251986 338614
rect 252222 338378 252306 338614
rect 252542 338378 271986 338614
rect 272222 338378 272306 338614
rect 272542 338378 291986 338614
rect 292222 338378 292306 338614
rect 292542 338378 311986 338614
rect 312222 338378 312306 338614
rect 312542 338378 331986 338614
rect 332222 338378 332306 338614
rect 332542 338378 351986 338614
rect 352222 338378 352306 338614
rect 352542 338378 371986 338614
rect 372222 338378 372306 338614
rect 372542 338378 391986 338614
rect 392222 338378 392306 338614
rect 392542 338378 411986 338614
rect 412222 338378 412306 338614
rect 412542 338378 431986 338614
rect 432222 338378 432306 338614
rect 432542 338378 451986 338614
rect 452222 338378 452306 338614
rect 452542 338378 471986 338614
rect 472222 338378 472306 338614
rect 472542 338378 491986 338614
rect 492222 338378 492306 338614
rect 492542 338378 511986 338614
rect 512222 338378 512306 338614
rect 512542 338378 531986 338614
rect 532222 338378 532306 338614
rect 532542 338378 551986 338614
rect 552222 338378 552306 338614
rect 552542 338378 571986 338614
rect 572222 338378 572306 338614
rect 572542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 11986 338294
rect 12222 338058 12306 338294
rect 12542 338058 31986 338294
rect 32222 338058 32306 338294
rect 32542 338058 51986 338294
rect 52222 338058 52306 338294
rect 52542 338058 71986 338294
rect 72222 338058 72306 338294
rect 72542 338058 91986 338294
rect 92222 338058 92306 338294
rect 92542 338058 111986 338294
rect 112222 338058 112306 338294
rect 112542 338058 131986 338294
rect 132222 338058 132306 338294
rect 132542 338058 151986 338294
rect 152222 338058 152306 338294
rect 152542 338058 171986 338294
rect 172222 338058 172306 338294
rect 172542 338058 191986 338294
rect 192222 338058 192306 338294
rect 192542 338058 211986 338294
rect 212222 338058 212306 338294
rect 212542 338058 231986 338294
rect 232222 338058 232306 338294
rect 232542 338058 251986 338294
rect 252222 338058 252306 338294
rect 252542 338058 271986 338294
rect 272222 338058 272306 338294
rect 272542 338058 291986 338294
rect 292222 338058 292306 338294
rect 292542 338058 311986 338294
rect 312222 338058 312306 338294
rect 312542 338058 331986 338294
rect 332222 338058 332306 338294
rect 332542 338058 351986 338294
rect 352222 338058 352306 338294
rect 352542 338058 371986 338294
rect 372222 338058 372306 338294
rect 372542 338058 391986 338294
rect 392222 338058 392306 338294
rect 392542 338058 411986 338294
rect 412222 338058 412306 338294
rect 412542 338058 431986 338294
rect 432222 338058 432306 338294
rect 432542 338058 451986 338294
rect 452222 338058 452306 338294
rect 452542 338058 471986 338294
rect 472222 338058 472306 338294
rect 472542 338058 491986 338294
rect 492222 338058 492306 338294
rect 492542 338058 511986 338294
rect 512222 338058 512306 338294
rect 512542 338058 531986 338294
rect 532222 338058 532306 338294
rect 532542 338058 551986 338294
rect 552222 338058 552306 338294
rect 552542 338058 571986 338294
rect 572222 338058 572306 338294
rect 572542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 8266 334894
rect 8502 334658 8586 334894
rect 8822 334658 28266 334894
rect 28502 334658 28586 334894
rect 28822 334658 48266 334894
rect 48502 334658 48586 334894
rect 48822 334658 68266 334894
rect 68502 334658 68586 334894
rect 68822 334658 88266 334894
rect 88502 334658 88586 334894
rect 88822 334658 108266 334894
rect 108502 334658 108586 334894
rect 108822 334658 128266 334894
rect 128502 334658 128586 334894
rect 128822 334658 148266 334894
rect 148502 334658 148586 334894
rect 148822 334658 168266 334894
rect 168502 334658 168586 334894
rect 168822 334658 188266 334894
rect 188502 334658 188586 334894
rect 188822 334658 208266 334894
rect 208502 334658 208586 334894
rect 208822 334658 228266 334894
rect 228502 334658 228586 334894
rect 228822 334658 248266 334894
rect 248502 334658 248586 334894
rect 248822 334658 268266 334894
rect 268502 334658 268586 334894
rect 268822 334658 288266 334894
rect 288502 334658 288586 334894
rect 288822 334658 308266 334894
rect 308502 334658 308586 334894
rect 308822 334658 328266 334894
rect 328502 334658 328586 334894
rect 328822 334658 348266 334894
rect 348502 334658 348586 334894
rect 348822 334658 368266 334894
rect 368502 334658 368586 334894
rect 368822 334658 388266 334894
rect 388502 334658 388586 334894
rect 388822 334658 408266 334894
rect 408502 334658 408586 334894
rect 408822 334658 428266 334894
rect 428502 334658 428586 334894
rect 428822 334658 448266 334894
rect 448502 334658 448586 334894
rect 448822 334658 468266 334894
rect 468502 334658 468586 334894
rect 468822 334658 488266 334894
rect 488502 334658 488586 334894
rect 488822 334658 508266 334894
rect 508502 334658 508586 334894
rect 508822 334658 528266 334894
rect 528502 334658 528586 334894
rect 528822 334658 548266 334894
rect 548502 334658 548586 334894
rect 548822 334658 568266 334894
rect 568502 334658 568586 334894
rect 568822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 8266 334574
rect 8502 334338 8586 334574
rect 8822 334338 28266 334574
rect 28502 334338 28586 334574
rect 28822 334338 48266 334574
rect 48502 334338 48586 334574
rect 48822 334338 68266 334574
rect 68502 334338 68586 334574
rect 68822 334338 88266 334574
rect 88502 334338 88586 334574
rect 88822 334338 108266 334574
rect 108502 334338 108586 334574
rect 108822 334338 128266 334574
rect 128502 334338 128586 334574
rect 128822 334338 148266 334574
rect 148502 334338 148586 334574
rect 148822 334338 168266 334574
rect 168502 334338 168586 334574
rect 168822 334338 188266 334574
rect 188502 334338 188586 334574
rect 188822 334338 208266 334574
rect 208502 334338 208586 334574
rect 208822 334338 228266 334574
rect 228502 334338 228586 334574
rect 228822 334338 248266 334574
rect 248502 334338 248586 334574
rect 248822 334338 268266 334574
rect 268502 334338 268586 334574
rect 268822 334338 288266 334574
rect 288502 334338 288586 334574
rect 288822 334338 308266 334574
rect 308502 334338 308586 334574
rect 308822 334338 328266 334574
rect 328502 334338 328586 334574
rect 328822 334338 348266 334574
rect 348502 334338 348586 334574
rect 348822 334338 368266 334574
rect 368502 334338 368586 334574
rect 368822 334338 388266 334574
rect 388502 334338 388586 334574
rect 388822 334338 408266 334574
rect 408502 334338 408586 334574
rect 408822 334338 428266 334574
rect 428502 334338 428586 334574
rect 428822 334338 448266 334574
rect 448502 334338 448586 334574
rect 448822 334338 468266 334574
rect 468502 334338 468586 334574
rect 468822 334338 488266 334574
rect 488502 334338 488586 334574
rect 488822 334338 508266 334574
rect 508502 334338 508586 334574
rect 508822 334338 528266 334574
rect 528502 334338 528586 334574
rect 528822 334338 548266 334574
rect 548502 334338 548586 334574
rect 548822 334338 568266 334574
rect 568502 334338 568586 334574
rect 568822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 4546 331174
rect 4782 330938 4866 331174
rect 5102 330938 24546 331174
rect 24782 330938 24866 331174
rect 25102 330938 44546 331174
rect 44782 330938 44866 331174
rect 45102 330938 64546 331174
rect 64782 330938 64866 331174
rect 65102 330938 84546 331174
rect 84782 330938 84866 331174
rect 85102 330938 104546 331174
rect 104782 330938 104866 331174
rect 105102 330938 124546 331174
rect 124782 330938 124866 331174
rect 125102 330938 144546 331174
rect 144782 330938 144866 331174
rect 145102 330938 164546 331174
rect 164782 330938 164866 331174
rect 165102 330938 184546 331174
rect 184782 330938 184866 331174
rect 185102 330938 204546 331174
rect 204782 330938 204866 331174
rect 205102 330938 224546 331174
rect 224782 330938 224866 331174
rect 225102 330938 244546 331174
rect 244782 330938 244866 331174
rect 245102 330938 264546 331174
rect 264782 330938 264866 331174
rect 265102 330938 284546 331174
rect 284782 330938 284866 331174
rect 285102 330938 304546 331174
rect 304782 330938 304866 331174
rect 305102 330938 324546 331174
rect 324782 330938 324866 331174
rect 325102 330938 344546 331174
rect 344782 330938 344866 331174
rect 345102 330938 364546 331174
rect 364782 330938 364866 331174
rect 365102 330938 384546 331174
rect 384782 330938 384866 331174
rect 385102 330938 404546 331174
rect 404782 330938 404866 331174
rect 405102 330938 424546 331174
rect 424782 330938 424866 331174
rect 425102 330938 444546 331174
rect 444782 330938 444866 331174
rect 445102 330938 464546 331174
rect 464782 330938 464866 331174
rect 465102 330938 484546 331174
rect 484782 330938 484866 331174
rect 485102 330938 504546 331174
rect 504782 330938 504866 331174
rect 505102 330938 524546 331174
rect 524782 330938 524866 331174
rect 525102 330938 544546 331174
rect 544782 330938 544866 331174
rect 545102 330938 564546 331174
rect 564782 330938 564866 331174
rect 565102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 4546 330854
rect 4782 330618 4866 330854
rect 5102 330618 24546 330854
rect 24782 330618 24866 330854
rect 25102 330618 44546 330854
rect 44782 330618 44866 330854
rect 45102 330618 64546 330854
rect 64782 330618 64866 330854
rect 65102 330618 84546 330854
rect 84782 330618 84866 330854
rect 85102 330618 104546 330854
rect 104782 330618 104866 330854
rect 105102 330618 124546 330854
rect 124782 330618 124866 330854
rect 125102 330618 144546 330854
rect 144782 330618 144866 330854
rect 145102 330618 164546 330854
rect 164782 330618 164866 330854
rect 165102 330618 184546 330854
rect 184782 330618 184866 330854
rect 185102 330618 204546 330854
rect 204782 330618 204866 330854
rect 205102 330618 224546 330854
rect 224782 330618 224866 330854
rect 225102 330618 244546 330854
rect 244782 330618 244866 330854
rect 245102 330618 264546 330854
rect 264782 330618 264866 330854
rect 265102 330618 284546 330854
rect 284782 330618 284866 330854
rect 285102 330618 304546 330854
rect 304782 330618 304866 330854
rect 305102 330618 324546 330854
rect 324782 330618 324866 330854
rect 325102 330618 344546 330854
rect 344782 330618 344866 330854
rect 345102 330618 364546 330854
rect 364782 330618 364866 330854
rect 365102 330618 384546 330854
rect 384782 330618 384866 330854
rect 385102 330618 404546 330854
rect 404782 330618 404866 330854
rect 405102 330618 424546 330854
rect 424782 330618 424866 330854
rect 425102 330618 444546 330854
rect 444782 330618 444866 330854
rect 445102 330618 464546 330854
rect 464782 330618 464866 330854
rect 465102 330618 484546 330854
rect 484782 330618 484866 330854
rect 485102 330618 504546 330854
rect 504782 330618 504866 330854
rect 505102 330618 524546 330854
rect 524782 330618 524866 330854
rect 525102 330618 544546 330854
rect 544782 330618 544866 330854
rect 545102 330618 564546 330854
rect 564782 330618 564866 330854
rect 565102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 826 327454
rect 1062 327218 1146 327454
rect 1382 327218 20826 327454
rect 21062 327218 21146 327454
rect 21382 327218 40826 327454
rect 41062 327218 41146 327454
rect 41382 327218 60826 327454
rect 61062 327218 61146 327454
rect 61382 327218 80826 327454
rect 81062 327218 81146 327454
rect 81382 327218 100826 327454
rect 101062 327218 101146 327454
rect 101382 327218 120826 327454
rect 121062 327218 121146 327454
rect 121382 327218 140826 327454
rect 141062 327218 141146 327454
rect 141382 327218 160826 327454
rect 161062 327218 161146 327454
rect 161382 327218 180826 327454
rect 181062 327218 181146 327454
rect 181382 327218 200826 327454
rect 201062 327218 201146 327454
rect 201382 327218 220826 327454
rect 221062 327218 221146 327454
rect 221382 327218 240826 327454
rect 241062 327218 241146 327454
rect 241382 327218 260826 327454
rect 261062 327218 261146 327454
rect 261382 327218 280826 327454
rect 281062 327218 281146 327454
rect 281382 327218 300826 327454
rect 301062 327218 301146 327454
rect 301382 327218 320826 327454
rect 321062 327218 321146 327454
rect 321382 327218 340826 327454
rect 341062 327218 341146 327454
rect 341382 327218 360826 327454
rect 361062 327218 361146 327454
rect 361382 327218 380826 327454
rect 381062 327218 381146 327454
rect 381382 327218 400826 327454
rect 401062 327218 401146 327454
rect 401382 327218 420826 327454
rect 421062 327218 421146 327454
rect 421382 327218 440826 327454
rect 441062 327218 441146 327454
rect 441382 327218 460826 327454
rect 461062 327218 461146 327454
rect 461382 327218 480826 327454
rect 481062 327218 481146 327454
rect 481382 327218 500826 327454
rect 501062 327218 501146 327454
rect 501382 327218 520826 327454
rect 521062 327218 521146 327454
rect 521382 327218 540826 327454
rect 541062 327218 541146 327454
rect 541382 327218 560826 327454
rect 561062 327218 561146 327454
rect 561382 327218 580826 327454
rect 581062 327218 581146 327454
rect 581382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 826 327134
rect 1062 326898 1146 327134
rect 1382 326898 20826 327134
rect 21062 326898 21146 327134
rect 21382 326898 40826 327134
rect 41062 326898 41146 327134
rect 41382 326898 60826 327134
rect 61062 326898 61146 327134
rect 61382 326898 80826 327134
rect 81062 326898 81146 327134
rect 81382 326898 100826 327134
rect 101062 326898 101146 327134
rect 101382 326898 120826 327134
rect 121062 326898 121146 327134
rect 121382 326898 140826 327134
rect 141062 326898 141146 327134
rect 141382 326898 160826 327134
rect 161062 326898 161146 327134
rect 161382 326898 180826 327134
rect 181062 326898 181146 327134
rect 181382 326898 200826 327134
rect 201062 326898 201146 327134
rect 201382 326898 220826 327134
rect 221062 326898 221146 327134
rect 221382 326898 240826 327134
rect 241062 326898 241146 327134
rect 241382 326898 260826 327134
rect 261062 326898 261146 327134
rect 261382 326898 280826 327134
rect 281062 326898 281146 327134
rect 281382 326898 300826 327134
rect 301062 326898 301146 327134
rect 301382 326898 320826 327134
rect 321062 326898 321146 327134
rect 321382 326898 340826 327134
rect 341062 326898 341146 327134
rect 341382 326898 360826 327134
rect 361062 326898 361146 327134
rect 361382 326898 380826 327134
rect 381062 326898 381146 327134
rect 381382 326898 400826 327134
rect 401062 326898 401146 327134
rect 401382 326898 420826 327134
rect 421062 326898 421146 327134
rect 421382 326898 440826 327134
rect 441062 326898 441146 327134
rect 441382 326898 460826 327134
rect 461062 326898 461146 327134
rect 461382 326898 480826 327134
rect 481062 326898 481146 327134
rect 481382 326898 500826 327134
rect 501062 326898 501146 327134
rect 501382 326898 520826 327134
rect 521062 326898 521146 327134
rect 521382 326898 540826 327134
rect 541062 326898 541146 327134
rect 541382 326898 560826 327134
rect 561062 326898 561146 327134
rect 561382 326898 580826 327134
rect 581062 326898 581146 327134
rect 581382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 21986 320614
rect 22222 320378 22306 320614
rect 22542 320378 41986 320614
rect 42222 320378 42306 320614
rect 42542 320378 61986 320614
rect 62222 320378 62306 320614
rect 62542 320378 81986 320614
rect 82222 320378 82306 320614
rect 82542 320378 101986 320614
rect 102222 320378 102306 320614
rect 102542 320378 121986 320614
rect 122222 320378 122306 320614
rect 122542 320378 141986 320614
rect 142222 320378 142306 320614
rect 142542 320378 161986 320614
rect 162222 320378 162306 320614
rect 162542 320378 181986 320614
rect 182222 320378 182306 320614
rect 182542 320378 201986 320614
rect 202222 320378 202306 320614
rect 202542 320378 221986 320614
rect 222222 320378 222306 320614
rect 222542 320378 241986 320614
rect 242222 320378 242306 320614
rect 242542 320378 261986 320614
rect 262222 320378 262306 320614
rect 262542 320378 281986 320614
rect 282222 320378 282306 320614
rect 282542 320378 301986 320614
rect 302222 320378 302306 320614
rect 302542 320378 321986 320614
rect 322222 320378 322306 320614
rect 322542 320378 341986 320614
rect 342222 320378 342306 320614
rect 342542 320378 361986 320614
rect 362222 320378 362306 320614
rect 362542 320378 381986 320614
rect 382222 320378 382306 320614
rect 382542 320378 401986 320614
rect 402222 320378 402306 320614
rect 402542 320378 421986 320614
rect 422222 320378 422306 320614
rect 422542 320378 441986 320614
rect 442222 320378 442306 320614
rect 442542 320378 461986 320614
rect 462222 320378 462306 320614
rect 462542 320378 481986 320614
rect 482222 320378 482306 320614
rect 482542 320378 501986 320614
rect 502222 320378 502306 320614
rect 502542 320378 521986 320614
rect 522222 320378 522306 320614
rect 522542 320378 541986 320614
rect 542222 320378 542306 320614
rect 542542 320378 561986 320614
rect 562222 320378 562306 320614
rect 562542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 21986 320294
rect 22222 320058 22306 320294
rect 22542 320058 41986 320294
rect 42222 320058 42306 320294
rect 42542 320058 61986 320294
rect 62222 320058 62306 320294
rect 62542 320058 81986 320294
rect 82222 320058 82306 320294
rect 82542 320058 101986 320294
rect 102222 320058 102306 320294
rect 102542 320058 121986 320294
rect 122222 320058 122306 320294
rect 122542 320058 141986 320294
rect 142222 320058 142306 320294
rect 142542 320058 161986 320294
rect 162222 320058 162306 320294
rect 162542 320058 181986 320294
rect 182222 320058 182306 320294
rect 182542 320058 201986 320294
rect 202222 320058 202306 320294
rect 202542 320058 221986 320294
rect 222222 320058 222306 320294
rect 222542 320058 241986 320294
rect 242222 320058 242306 320294
rect 242542 320058 261986 320294
rect 262222 320058 262306 320294
rect 262542 320058 281986 320294
rect 282222 320058 282306 320294
rect 282542 320058 301986 320294
rect 302222 320058 302306 320294
rect 302542 320058 321986 320294
rect 322222 320058 322306 320294
rect 322542 320058 341986 320294
rect 342222 320058 342306 320294
rect 342542 320058 361986 320294
rect 362222 320058 362306 320294
rect 362542 320058 381986 320294
rect 382222 320058 382306 320294
rect 382542 320058 401986 320294
rect 402222 320058 402306 320294
rect 402542 320058 421986 320294
rect 422222 320058 422306 320294
rect 422542 320058 441986 320294
rect 442222 320058 442306 320294
rect 442542 320058 461986 320294
rect 462222 320058 462306 320294
rect 462542 320058 481986 320294
rect 482222 320058 482306 320294
rect 482542 320058 501986 320294
rect 502222 320058 502306 320294
rect 502542 320058 521986 320294
rect 522222 320058 522306 320294
rect 522542 320058 541986 320294
rect 542222 320058 542306 320294
rect 542542 320058 561986 320294
rect 562222 320058 562306 320294
rect 562542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 18266 316894
rect 18502 316658 18586 316894
rect 18822 316658 38266 316894
rect 38502 316658 38586 316894
rect 38822 316658 58266 316894
rect 58502 316658 58586 316894
rect 58822 316658 78266 316894
rect 78502 316658 78586 316894
rect 78822 316658 98266 316894
rect 98502 316658 98586 316894
rect 98822 316658 118266 316894
rect 118502 316658 118586 316894
rect 118822 316658 138266 316894
rect 138502 316658 138586 316894
rect 138822 316658 158266 316894
rect 158502 316658 158586 316894
rect 158822 316658 178266 316894
rect 178502 316658 178586 316894
rect 178822 316658 198266 316894
rect 198502 316658 198586 316894
rect 198822 316658 218266 316894
rect 218502 316658 218586 316894
rect 218822 316658 238266 316894
rect 238502 316658 238586 316894
rect 238822 316658 258266 316894
rect 258502 316658 258586 316894
rect 258822 316658 278266 316894
rect 278502 316658 278586 316894
rect 278822 316658 298266 316894
rect 298502 316658 298586 316894
rect 298822 316658 318266 316894
rect 318502 316658 318586 316894
rect 318822 316658 338266 316894
rect 338502 316658 338586 316894
rect 338822 316658 358266 316894
rect 358502 316658 358586 316894
rect 358822 316658 378266 316894
rect 378502 316658 378586 316894
rect 378822 316658 398266 316894
rect 398502 316658 398586 316894
rect 398822 316658 418266 316894
rect 418502 316658 418586 316894
rect 418822 316658 438266 316894
rect 438502 316658 438586 316894
rect 438822 316658 458266 316894
rect 458502 316658 458586 316894
rect 458822 316658 478266 316894
rect 478502 316658 478586 316894
rect 478822 316658 498266 316894
rect 498502 316658 498586 316894
rect 498822 316658 518266 316894
rect 518502 316658 518586 316894
rect 518822 316658 538266 316894
rect 538502 316658 538586 316894
rect 538822 316658 558266 316894
rect 558502 316658 558586 316894
rect 558822 316658 578266 316894
rect 578502 316658 578586 316894
rect 578822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 18266 316574
rect 18502 316338 18586 316574
rect 18822 316338 38266 316574
rect 38502 316338 38586 316574
rect 38822 316338 58266 316574
rect 58502 316338 58586 316574
rect 58822 316338 78266 316574
rect 78502 316338 78586 316574
rect 78822 316338 98266 316574
rect 98502 316338 98586 316574
rect 98822 316338 118266 316574
rect 118502 316338 118586 316574
rect 118822 316338 138266 316574
rect 138502 316338 138586 316574
rect 138822 316338 158266 316574
rect 158502 316338 158586 316574
rect 158822 316338 178266 316574
rect 178502 316338 178586 316574
rect 178822 316338 198266 316574
rect 198502 316338 198586 316574
rect 198822 316338 218266 316574
rect 218502 316338 218586 316574
rect 218822 316338 238266 316574
rect 238502 316338 238586 316574
rect 238822 316338 258266 316574
rect 258502 316338 258586 316574
rect 258822 316338 278266 316574
rect 278502 316338 278586 316574
rect 278822 316338 298266 316574
rect 298502 316338 298586 316574
rect 298822 316338 318266 316574
rect 318502 316338 318586 316574
rect 318822 316338 338266 316574
rect 338502 316338 338586 316574
rect 338822 316338 358266 316574
rect 358502 316338 358586 316574
rect 358822 316338 378266 316574
rect 378502 316338 378586 316574
rect 378822 316338 398266 316574
rect 398502 316338 398586 316574
rect 398822 316338 418266 316574
rect 418502 316338 418586 316574
rect 418822 316338 438266 316574
rect 438502 316338 438586 316574
rect 438822 316338 458266 316574
rect 458502 316338 458586 316574
rect 458822 316338 478266 316574
rect 478502 316338 478586 316574
rect 478822 316338 498266 316574
rect 498502 316338 498586 316574
rect 498822 316338 518266 316574
rect 518502 316338 518586 316574
rect 518822 316338 538266 316574
rect 538502 316338 538586 316574
rect 538822 316338 558266 316574
rect 558502 316338 558586 316574
rect 558822 316338 578266 316574
rect 578502 316338 578586 316574
rect 578822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 14546 313174
rect 14782 312938 14866 313174
rect 15102 312938 34546 313174
rect 34782 312938 34866 313174
rect 35102 312938 54546 313174
rect 54782 312938 54866 313174
rect 55102 312938 74546 313174
rect 74782 312938 74866 313174
rect 75102 312938 94546 313174
rect 94782 312938 94866 313174
rect 95102 312938 114546 313174
rect 114782 312938 114866 313174
rect 115102 312938 134546 313174
rect 134782 312938 134866 313174
rect 135102 312938 154546 313174
rect 154782 312938 154866 313174
rect 155102 312938 174546 313174
rect 174782 312938 174866 313174
rect 175102 312938 194546 313174
rect 194782 312938 194866 313174
rect 195102 312938 214546 313174
rect 214782 312938 214866 313174
rect 215102 312938 234546 313174
rect 234782 312938 234866 313174
rect 235102 312938 254546 313174
rect 254782 312938 254866 313174
rect 255102 312938 274546 313174
rect 274782 312938 274866 313174
rect 275102 312938 294546 313174
rect 294782 312938 294866 313174
rect 295102 312938 314546 313174
rect 314782 312938 314866 313174
rect 315102 312938 334546 313174
rect 334782 312938 334866 313174
rect 335102 312938 354546 313174
rect 354782 312938 354866 313174
rect 355102 312938 374546 313174
rect 374782 312938 374866 313174
rect 375102 312938 394546 313174
rect 394782 312938 394866 313174
rect 395102 312938 414546 313174
rect 414782 312938 414866 313174
rect 415102 312938 434546 313174
rect 434782 312938 434866 313174
rect 435102 312938 454546 313174
rect 454782 312938 454866 313174
rect 455102 312938 474546 313174
rect 474782 312938 474866 313174
rect 475102 312938 494546 313174
rect 494782 312938 494866 313174
rect 495102 312938 514546 313174
rect 514782 312938 514866 313174
rect 515102 312938 534546 313174
rect 534782 312938 534866 313174
rect 535102 312938 554546 313174
rect 554782 312938 554866 313174
rect 555102 312938 574546 313174
rect 574782 312938 574866 313174
rect 575102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 14546 312854
rect 14782 312618 14866 312854
rect 15102 312618 34546 312854
rect 34782 312618 34866 312854
rect 35102 312618 54546 312854
rect 54782 312618 54866 312854
rect 55102 312618 74546 312854
rect 74782 312618 74866 312854
rect 75102 312618 94546 312854
rect 94782 312618 94866 312854
rect 95102 312618 114546 312854
rect 114782 312618 114866 312854
rect 115102 312618 134546 312854
rect 134782 312618 134866 312854
rect 135102 312618 154546 312854
rect 154782 312618 154866 312854
rect 155102 312618 174546 312854
rect 174782 312618 174866 312854
rect 175102 312618 194546 312854
rect 194782 312618 194866 312854
rect 195102 312618 214546 312854
rect 214782 312618 214866 312854
rect 215102 312618 234546 312854
rect 234782 312618 234866 312854
rect 235102 312618 254546 312854
rect 254782 312618 254866 312854
rect 255102 312618 274546 312854
rect 274782 312618 274866 312854
rect 275102 312618 294546 312854
rect 294782 312618 294866 312854
rect 295102 312618 314546 312854
rect 314782 312618 314866 312854
rect 315102 312618 334546 312854
rect 334782 312618 334866 312854
rect 335102 312618 354546 312854
rect 354782 312618 354866 312854
rect 355102 312618 374546 312854
rect 374782 312618 374866 312854
rect 375102 312618 394546 312854
rect 394782 312618 394866 312854
rect 395102 312618 414546 312854
rect 414782 312618 414866 312854
rect 415102 312618 434546 312854
rect 434782 312618 434866 312854
rect 435102 312618 454546 312854
rect 454782 312618 454866 312854
rect 455102 312618 474546 312854
rect 474782 312618 474866 312854
rect 475102 312618 494546 312854
rect 494782 312618 494866 312854
rect 495102 312618 514546 312854
rect 514782 312618 514866 312854
rect 515102 312618 534546 312854
rect 534782 312618 534866 312854
rect 535102 312618 554546 312854
rect 554782 312618 554866 312854
rect 555102 312618 574546 312854
rect 574782 312618 574866 312854
rect 575102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 10826 309454
rect 11062 309218 11146 309454
rect 11382 309218 30826 309454
rect 31062 309218 31146 309454
rect 31382 309218 50826 309454
rect 51062 309218 51146 309454
rect 51382 309218 70826 309454
rect 71062 309218 71146 309454
rect 71382 309218 90826 309454
rect 91062 309218 91146 309454
rect 91382 309218 110826 309454
rect 111062 309218 111146 309454
rect 111382 309218 130826 309454
rect 131062 309218 131146 309454
rect 131382 309218 150826 309454
rect 151062 309218 151146 309454
rect 151382 309218 170826 309454
rect 171062 309218 171146 309454
rect 171382 309218 190826 309454
rect 191062 309218 191146 309454
rect 191382 309218 210826 309454
rect 211062 309218 211146 309454
rect 211382 309218 230826 309454
rect 231062 309218 231146 309454
rect 231382 309218 250826 309454
rect 251062 309218 251146 309454
rect 251382 309218 270826 309454
rect 271062 309218 271146 309454
rect 271382 309218 290826 309454
rect 291062 309218 291146 309454
rect 291382 309218 310826 309454
rect 311062 309218 311146 309454
rect 311382 309218 330826 309454
rect 331062 309218 331146 309454
rect 331382 309218 350826 309454
rect 351062 309218 351146 309454
rect 351382 309218 370826 309454
rect 371062 309218 371146 309454
rect 371382 309218 390826 309454
rect 391062 309218 391146 309454
rect 391382 309218 410826 309454
rect 411062 309218 411146 309454
rect 411382 309218 430826 309454
rect 431062 309218 431146 309454
rect 431382 309218 450826 309454
rect 451062 309218 451146 309454
rect 451382 309218 470826 309454
rect 471062 309218 471146 309454
rect 471382 309218 490826 309454
rect 491062 309218 491146 309454
rect 491382 309218 510826 309454
rect 511062 309218 511146 309454
rect 511382 309218 530826 309454
rect 531062 309218 531146 309454
rect 531382 309218 550826 309454
rect 551062 309218 551146 309454
rect 551382 309218 570826 309454
rect 571062 309218 571146 309454
rect 571382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 10826 309134
rect 11062 308898 11146 309134
rect 11382 308898 30826 309134
rect 31062 308898 31146 309134
rect 31382 308898 50826 309134
rect 51062 308898 51146 309134
rect 51382 308898 70826 309134
rect 71062 308898 71146 309134
rect 71382 308898 90826 309134
rect 91062 308898 91146 309134
rect 91382 308898 110826 309134
rect 111062 308898 111146 309134
rect 111382 308898 130826 309134
rect 131062 308898 131146 309134
rect 131382 308898 150826 309134
rect 151062 308898 151146 309134
rect 151382 308898 170826 309134
rect 171062 308898 171146 309134
rect 171382 308898 190826 309134
rect 191062 308898 191146 309134
rect 191382 308898 210826 309134
rect 211062 308898 211146 309134
rect 211382 308898 230826 309134
rect 231062 308898 231146 309134
rect 231382 308898 250826 309134
rect 251062 308898 251146 309134
rect 251382 308898 270826 309134
rect 271062 308898 271146 309134
rect 271382 308898 290826 309134
rect 291062 308898 291146 309134
rect 291382 308898 310826 309134
rect 311062 308898 311146 309134
rect 311382 308898 330826 309134
rect 331062 308898 331146 309134
rect 331382 308898 350826 309134
rect 351062 308898 351146 309134
rect 351382 308898 370826 309134
rect 371062 308898 371146 309134
rect 371382 308898 390826 309134
rect 391062 308898 391146 309134
rect 391382 308898 410826 309134
rect 411062 308898 411146 309134
rect 411382 308898 430826 309134
rect 431062 308898 431146 309134
rect 431382 308898 450826 309134
rect 451062 308898 451146 309134
rect 451382 308898 470826 309134
rect 471062 308898 471146 309134
rect 471382 308898 490826 309134
rect 491062 308898 491146 309134
rect 491382 308898 510826 309134
rect 511062 308898 511146 309134
rect 511382 308898 530826 309134
rect 531062 308898 531146 309134
rect 531382 308898 550826 309134
rect 551062 308898 551146 309134
rect 551382 308898 570826 309134
rect 571062 308898 571146 309134
rect 571382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 11986 302614
rect 12222 302378 12306 302614
rect 12542 302378 31986 302614
rect 32222 302378 32306 302614
rect 32542 302378 51986 302614
rect 52222 302378 52306 302614
rect 52542 302378 71986 302614
rect 72222 302378 72306 302614
rect 72542 302378 91986 302614
rect 92222 302378 92306 302614
rect 92542 302378 111986 302614
rect 112222 302378 112306 302614
rect 112542 302378 131986 302614
rect 132222 302378 132306 302614
rect 132542 302378 151986 302614
rect 152222 302378 152306 302614
rect 152542 302378 171986 302614
rect 172222 302378 172306 302614
rect 172542 302378 191986 302614
rect 192222 302378 192306 302614
rect 192542 302378 211986 302614
rect 212222 302378 212306 302614
rect 212542 302378 231986 302614
rect 232222 302378 232306 302614
rect 232542 302378 251986 302614
rect 252222 302378 252306 302614
rect 252542 302378 271986 302614
rect 272222 302378 272306 302614
rect 272542 302378 291986 302614
rect 292222 302378 292306 302614
rect 292542 302378 311986 302614
rect 312222 302378 312306 302614
rect 312542 302378 331986 302614
rect 332222 302378 332306 302614
rect 332542 302378 351986 302614
rect 352222 302378 352306 302614
rect 352542 302378 371986 302614
rect 372222 302378 372306 302614
rect 372542 302378 391986 302614
rect 392222 302378 392306 302614
rect 392542 302378 411986 302614
rect 412222 302378 412306 302614
rect 412542 302378 431986 302614
rect 432222 302378 432306 302614
rect 432542 302378 451986 302614
rect 452222 302378 452306 302614
rect 452542 302378 471986 302614
rect 472222 302378 472306 302614
rect 472542 302378 491986 302614
rect 492222 302378 492306 302614
rect 492542 302378 511986 302614
rect 512222 302378 512306 302614
rect 512542 302378 531986 302614
rect 532222 302378 532306 302614
rect 532542 302378 551986 302614
rect 552222 302378 552306 302614
rect 552542 302378 571986 302614
rect 572222 302378 572306 302614
rect 572542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 11986 302294
rect 12222 302058 12306 302294
rect 12542 302058 31986 302294
rect 32222 302058 32306 302294
rect 32542 302058 51986 302294
rect 52222 302058 52306 302294
rect 52542 302058 71986 302294
rect 72222 302058 72306 302294
rect 72542 302058 91986 302294
rect 92222 302058 92306 302294
rect 92542 302058 111986 302294
rect 112222 302058 112306 302294
rect 112542 302058 131986 302294
rect 132222 302058 132306 302294
rect 132542 302058 151986 302294
rect 152222 302058 152306 302294
rect 152542 302058 171986 302294
rect 172222 302058 172306 302294
rect 172542 302058 191986 302294
rect 192222 302058 192306 302294
rect 192542 302058 211986 302294
rect 212222 302058 212306 302294
rect 212542 302058 231986 302294
rect 232222 302058 232306 302294
rect 232542 302058 251986 302294
rect 252222 302058 252306 302294
rect 252542 302058 271986 302294
rect 272222 302058 272306 302294
rect 272542 302058 291986 302294
rect 292222 302058 292306 302294
rect 292542 302058 311986 302294
rect 312222 302058 312306 302294
rect 312542 302058 331986 302294
rect 332222 302058 332306 302294
rect 332542 302058 351986 302294
rect 352222 302058 352306 302294
rect 352542 302058 371986 302294
rect 372222 302058 372306 302294
rect 372542 302058 391986 302294
rect 392222 302058 392306 302294
rect 392542 302058 411986 302294
rect 412222 302058 412306 302294
rect 412542 302058 431986 302294
rect 432222 302058 432306 302294
rect 432542 302058 451986 302294
rect 452222 302058 452306 302294
rect 452542 302058 471986 302294
rect 472222 302058 472306 302294
rect 472542 302058 491986 302294
rect 492222 302058 492306 302294
rect 492542 302058 511986 302294
rect 512222 302058 512306 302294
rect 512542 302058 531986 302294
rect 532222 302058 532306 302294
rect 532542 302058 551986 302294
rect 552222 302058 552306 302294
rect 552542 302058 571986 302294
rect 572222 302058 572306 302294
rect 572542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 8266 298894
rect 8502 298658 8586 298894
rect 8822 298658 28266 298894
rect 28502 298658 28586 298894
rect 28822 298658 48266 298894
rect 48502 298658 48586 298894
rect 48822 298658 68266 298894
rect 68502 298658 68586 298894
rect 68822 298658 88266 298894
rect 88502 298658 88586 298894
rect 88822 298658 108266 298894
rect 108502 298658 108586 298894
rect 108822 298658 128266 298894
rect 128502 298658 128586 298894
rect 128822 298658 148266 298894
rect 148502 298658 148586 298894
rect 148822 298658 168266 298894
rect 168502 298658 168586 298894
rect 168822 298658 188266 298894
rect 188502 298658 188586 298894
rect 188822 298658 208266 298894
rect 208502 298658 208586 298894
rect 208822 298658 228266 298894
rect 228502 298658 228586 298894
rect 228822 298658 248266 298894
rect 248502 298658 248586 298894
rect 248822 298658 268266 298894
rect 268502 298658 268586 298894
rect 268822 298658 288266 298894
rect 288502 298658 288586 298894
rect 288822 298658 308266 298894
rect 308502 298658 308586 298894
rect 308822 298658 328266 298894
rect 328502 298658 328586 298894
rect 328822 298658 348266 298894
rect 348502 298658 348586 298894
rect 348822 298658 368266 298894
rect 368502 298658 368586 298894
rect 368822 298658 388266 298894
rect 388502 298658 388586 298894
rect 388822 298658 408266 298894
rect 408502 298658 408586 298894
rect 408822 298658 428266 298894
rect 428502 298658 428586 298894
rect 428822 298658 448266 298894
rect 448502 298658 448586 298894
rect 448822 298658 468266 298894
rect 468502 298658 468586 298894
rect 468822 298658 488266 298894
rect 488502 298658 488586 298894
rect 488822 298658 508266 298894
rect 508502 298658 508586 298894
rect 508822 298658 528266 298894
rect 528502 298658 528586 298894
rect 528822 298658 548266 298894
rect 548502 298658 548586 298894
rect 548822 298658 568266 298894
rect 568502 298658 568586 298894
rect 568822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 8266 298574
rect 8502 298338 8586 298574
rect 8822 298338 28266 298574
rect 28502 298338 28586 298574
rect 28822 298338 48266 298574
rect 48502 298338 48586 298574
rect 48822 298338 68266 298574
rect 68502 298338 68586 298574
rect 68822 298338 88266 298574
rect 88502 298338 88586 298574
rect 88822 298338 108266 298574
rect 108502 298338 108586 298574
rect 108822 298338 128266 298574
rect 128502 298338 128586 298574
rect 128822 298338 148266 298574
rect 148502 298338 148586 298574
rect 148822 298338 168266 298574
rect 168502 298338 168586 298574
rect 168822 298338 188266 298574
rect 188502 298338 188586 298574
rect 188822 298338 208266 298574
rect 208502 298338 208586 298574
rect 208822 298338 228266 298574
rect 228502 298338 228586 298574
rect 228822 298338 248266 298574
rect 248502 298338 248586 298574
rect 248822 298338 268266 298574
rect 268502 298338 268586 298574
rect 268822 298338 288266 298574
rect 288502 298338 288586 298574
rect 288822 298338 308266 298574
rect 308502 298338 308586 298574
rect 308822 298338 328266 298574
rect 328502 298338 328586 298574
rect 328822 298338 348266 298574
rect 348502 298338 348586 298574
rect 348822 298338 368266 298574
rect 368502 298338 368586 298574
rect 368822 298338 388266 298574
rect 388502 298338 388586 298574
rect 388822 298338 408266 298574
rect 408502 298338 408586 298574
rect 408822 298338 428266 298574
rect 428502 298338 428586 298574
rect 428822 298338 448266 298574
rect 448502 298338 448586 298574
rect 448822 298338 468266 298574
rect 468502 298338 468586 298574
rect 468822 298338 488266 298574
rect 488502 298338 488586 298574
rect 488822 298338 508266 298574
rect 508502 298338 508586 298574
rect 508822 298338 528266 298574
rect 528502 298338 528586 298574
rect 528822 298338 548266 298574
rect 548502 298338 548586 298574
rect 548822 298338 568266 298574
rect 568502 298338 568586 298574
rect 568822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 4546 295174
rect 4782 294938 4866 295174
rect 5102 294938 24546 295174
rect 24782 294938 24866 295174
rect 25102 294938 44546 295174
rect 44782 294938 44866 295174
rect 45102 294938 64546 295174
rect 64782 294938 64866 295174
rect 65102 294938 84546 295174
rect 84782 294938 84866 295174
rect 85102 294938 104546 295174
rect 104782 294938 104866 295174
rect 105102 294938 124546 295174
rect 124782 294938 124866 295174
rect 125102 294938 144546 295174
rect 144782 294938 144866 295174
rect 145102 294938 164546 295174
rect 164782 294938 164866 295174
rect 165102 294938 184546 295174
rect 184782 294938 184866 295174
rect 185102 294938 204546 295174
rect 204782 294938 204866 295174
rect 205102 294938 224546 295174
rect 224782 294938 224866 295174
rect 225102 294938 244546 295174
rect 244782 294938 244866 295174
rect 245102 294938 264546 295174
rect 264782 294938 264866 295174
rect 265102 294938 284546 295174
rect 284782 294938 284866 295174
rect 285102 294938 304546 295174
rect 304782 294938 304866 295174
rect 305102 294938 324546 295174
rect 324782 294938 324866 295174
rect 325102 294938 344546 295174
rect 344782 294938 344866 295174
rect 345102 294938 364546 295174
rect 364782 294938 364866 295174
rect 365102 294938 384546 295174
rect 384782 294938 384866 295174
rect 385102 294938 404546 295174
rect 404782 294938 404866 295174
rect 405102 294938 424546 295174
rect 424782 294938 424866 295174
rect 425102 294938 444546 295174
rect 444782 294938 444866 295174
rect 445102 294938 464546 295174
rect 464782 294938 464866 295174
rect 465102 294938 484546 295174
rect 484782 294938 484866 295174
rect 485102 294938 504546 295174
rect 504782 294938 504866 295174
rect 505102 294938 524546 295174
rect 524782 294938 524866 295174
rect 525102 294938 544546 295174
rect 544782 294938 544866 295174
rect 545102 294938 564546 295174
rect 564782 294938 564866 295174
rect 565102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 4546 294854
rect 4782 294618 4866 294854
rect 5102 294618 24546 294854
rect 24782 294618 24866 294854
rect 25102 294618 44546 294854
rect 44782 294618 44866 294854
rect 45102 294618 64546 294854
rect 64782 294618 64866 294854
rect 65102 294618 84546 294854
rect 84782 294618 84866 294854
rect 85102 294618 104546 294854
rect 104782 294618 104866 294854
rect 105102 294618 124546 294854
rect 124782 294618 124866 294854
rect 125102 294618 144546 294854
rect 144782 294618 144866 294854
rect 145102 294618 164546 294854
rect 164782 294618 164866 294854
rect 165102 294618 184546 294854
rect 184782 294618 184866 294854
rect 185102 294618 204546 294854
rect 204782 294618 204866 294854
rect 205102 294618 224546 294854
rect 224782 294618 224866 294854
rect 225102 294618 244546 294854
rect 244782 294618 244866 294854
rect 245102 294618 264546 294854
rect 264782 294618 264866 294854
rect 265102 294618 284546 294854
rect 284782 294618 284866 294854
rect 285102 294618 304546 294854
rect 304782 294618 304866 294854
rect 305102 294618 324546 294854
rect 324782 294618 324866 294854
rect 325102 294618 344546 294854
rect 344782 294618 344866 294854
rect 345102 294618 364546 294854
rect 364782 294618 364866 294854
rect 365102 294618 384546 294854
rect 384782 294618 384866 294854
rect 385102 294618 404546 294854
rect 404782 294618 404866 294854
rect 405102 294618 424546 294854
rect 424782 294618 424866 294854
rect 425102 294618 444546 294854
rect 444782 294618 444866 294854
rect 445102 294618 464546 294854
rect 464782 294618 464866 294854
rect 465102 294618 484546 294854
rect 484782 294618 484866 294854
rect 485102 294618 504546 294854
rect 504782 294618 504866 294854
rect 505102 294618 524546 294854
rect 524782 294618 524866 294854
rect 525102 294618 544546 294854
rect 544782 294618 544866 294854
rect 545102 294618 564546 294854
rect 564782 294618 564866 294854
rect 565102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 826 291454
rect 1062 291218 1146 291454
rect 1382 291218 20826 291454
rect 21062 291218 21146 291454
rect 21382 291218 40826 291454
rect 41062 291218 41146 291454
rect 41382 291218 60826 291454
rect 61062 291218 61146 291454
rect 61382 291218 80826 291454
rect 81062 291218 81146 291454
rect 81382 291218 100826 291454
rect 101062 291218 101146 291454
rect 101382 291218 120826 291454
rect 121062 291218 121146 291454
rect 121382 291218 140826 291454
rect 141062 291218 141146 291454
rect 141382 291218 160826 291454
rect 161062 291218 161146 291454
rect 161382 291218 180826 291454
rect 181062 291218 181146 291454
rect 181382 291218 200826 291454
rect 201062 291218 201146 291454
rect 201382 291218 220826 291454
rect 221062 291218 221146 291454
rect 221382 291218 240826 291454
rect 241062 291218 241146 291454
rect 241382 291218 260826 291454
rect 261062 291218 261146 291454
rect 261382 291218 280826 291454
rect 281062 291218 281146 291454
rect 281382 291218 300826 291454
rect 301062 291218 301146 291454
rect 301382 291218 320826 291454
rect 321062 291218 321146 291454
rect 321382 291218 340826 291454
rect 341062 291218 341146 291454
rect 341382 291218 360826 291454
rect 361062 291218 361146 291454
rect 361382 291218 380826 291454
rect 381062 291218 381146 291454
rect 381382 291218 400826 291454
rect 401062 291218 401146 291454
rect 401382 291218 420826 291454
rect 421062 291218 421146 291454
rect 421382 291218 440826 291454
rect 441062 291218 441146 291454
rect 441382 291218 460826 291454
rect 461062 291218 461146 291454
rect 461382 291218 480826 291454
rect 481062 291218 481146 291454
rect 481382 291218 500826 291454
rect 501062 291218 501146 291454
rect 501382 291218 520826 291454
rect 521062 291218 521146 291454
rect 521382 291218 540826 291454
rect 541062 291218 541146 291454
rect 541382 291218 560826 291454
rect 561062 291218 561146 291454
rect 561382 291218 580826 291454
rect 581062 291218 581146 291454
rect 581382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 826 291134
rect 1062 290898 1146 291134
rect 1382 290898 20826 291134
rect 21062 290898 21146 291134
rect 21382 290898 40826 291134
rect 41062 290898 41146 291134
rect 41382 290898 60826 291134
rect 61062 290898 61146 291134
rect 61382 290898 80826 291134
rect 81062 290898 81146 291134
rect 81382 290898 100826 291134
rect 101062 290898 101146 291134
rect 101382 290898 120826 291134
rect 121062 290898 121146 291134
rect 121382 290898 140826 291134
rect 141062 290898 141146 291134
rect 141382 290898 160826 291134
rect 161062 290898 161146 291134
rect 161382 290898 180826 291134
rect 181062 290898 181146 291134
rect 181382 290898 200826 291134
rect 201062 290898 201146 291134
rect 201382 290898 220826 291134
rect 221062 290898 221146 291134
rect 221382 290898 240826 291134
rect 241062 290898 241146 291134
rect 241382 290898 260826 291134
rect 261062 290898 261146 291134
rect 261382 290898 280826 291134
rect 281062 290898 281146 291134
rect 281382 290898 300826 291134
rect 301062 290898 301146 291134
rect 301382 290898 320826 291134
rect 321062 290898 321146 291134
rect 321382 290898 340826 291134
rect 341062 290898 341146 291134
rect 341382 290898 360826 291134
rect 361062 290898 361146 291134
rect 361382 290898 380826 291134
rect 381062 290898 381146 291134
rect 381382 290898 400826 291134
rect 401062 290898 401146 291134
rect 401382 290898 420826 291134
rect 421062 290898 421146 291134
rect 421382 290898 440826 291134
rect 441062 290898 441146 291134
rect 441382 290898 460826 291134
rect 461062 290898 461146 291134
rect 461382 290898 480826 291134
rect 481062 290898 481146 291134
rect 481382 290898 500826 291134
rect 501062 290898 501146 291134
rect 501382 290898 520826 291134
rect 521062 290898 521146 291134
rect 521382 290898 540826 291134
rect 541062 290898 541146 291134
rect 541382 290898 560826 291134
rect 561062 290898 561146 291134
rect 561382 290898 580826 291134
rect 581062 290898 581146 291134
rect 581382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 21986 284614
rect 22222 284378 22306 284614
rect 22542 284378 41986 284614
rect 42222 284378 42306 284614
rect 42542 284378 61986 284614
rect 62222 284378 62306 284614
rect 62542 284378 81986 284614
rect 82222 284378 82306 284614
rect 82542 284378 101986 284614
rect 102222 284378 102306 284614
rect 102542 284378 121986 284614
rect 122222 284378 122306 284614
rect 122542 284378 141986 284614
rect 142222 284378 142306 284614
rect 142542 284378 161986 284614
rect 162222 284378 162306 284614
rect 162542 284378 181986 284614
rect 182222 284378 182306 284614
rect 182542 284378 201986 284614
rect 202222 284378 202306 284614
rect 202542 284378 221986 284614
rect 222222 284378 222306 284614
rect 222542 284378 241986 284614
rect 242222 284378 242306 284614
rect 242542 284378 261986 284614
rect 262222 284378 262306 284614
rect 262542 284378 281986 284614
rect 282222 284378 282306 284614
rect 282542 284378 301986 284614
rect 302222 284378 302306 284614
rect 302542 284378 321986 284614
rect 322222 284378 322306 284614
rect 322542 284378 341986 284614
rect 342222 284378 342306 284614
rect 342542 284378 361986 284614
rect 362222 284378 362306 284614
rect 362542 284378 381986 284614
rect 382222 284378 382306 284614
rect 382542 284378 401986 284614
rect 402222 284378 402306 284614
rect 402542 284378 421986 284614
rect 422222 284378 422306 284614
rect 422542 284378 441986 284614
rect 442222 284378 442306 284614
rect 442542 284378 461986 284614
rect 462222 284378 462306 284614
rect 462542 284378 481986 284614
rect 482222 284378 482306 284614
rect 482542 284378 501986 284614
rect 502222 284378 502306 284614
rect 502542 284378 521986 284614
rect 522222 284378 522306 284614
rect 522542 284378 541986 284614
rect 542222 284378 542306 284614
rect 542542 284378 561986 284614
rect 562222 284378 562306 284614
rect 562542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 21986 284294
rect 22222 284058 22306 284294
rect 22542 284058 41986 284294
rect 42222 284058 42306 284294
rect 42542 284058 61986 284294
rect 62222 284058 62306 284294
rect 62542 284058 81986 284294
rect 82222 284058 82306 284294
rect 82542 284058 101986 284294
rect 102222 284058 102306 284294
rect 102542 284058 121986 284294
rect 122222 284058 122306 284294
rect 122542 284058 141986 284294
rect 142222 284058 142306 284294
rect 142542 284058 161986 284294
rect 162222 284058 162306 284294
rect 162542 284058 181986 284294
rect 182222 284058 182306 284294
rect 182542 284058 201986 284294
rect 202222 284058 202306 284294
rect 202542 284058 221986 284294
rect 222222 284058 222306 284294
rect 222542 284058 241986 284294
rect 242222 284058 242306 284294
rect 242542 284058 261986 284294
rect 262222 284058 262306 284294
rect 262542 284058 281986 284294
rect 282222 284058 282306 284294
rect 282542 284058 301986 284294
rect 302222 284058 302306 284294
rect 302542 284058 321986 284294
rect 322222 284058 322306 284294
rect 322542 284058 341986 284294
rect 342222 284058 342306 284294
rect 342542 284058 361986 284294
rect 362222 284058 362306 284294
rect 362542 284058 381986 284294
rect 382222 284058 382306 284294
rect 382542 284058 401986 284294
rect 402222 284058 402306 284294
rect 402542 284058 421986 284294
rect 422222 284058 422306 284294
rect 422542 284058 441986 284294
rect 442222 284058 442306 284294
rect 442542 284058 461986 284294
rect 462222 284058 462306 284294
rect 462542 284058 481986 284294
rect 482222 284058 482306 284294
rect 482542 284058 501986 284294
rect 502222 284058 502306 284294
rect 502542 284058 521986 284294
rect 522222 284058 522306 284294
rect 522542 284058 541986 284294
rect 542222 284058 542306 284294
rect 542542 284058 561986 284294
rect 562222 284058 562306 284294
rect 562542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 18266 280894
rect 18502 280658 18586 280894
rect 18822 280658 38266 280894
rect 38502 280658 38586 280894
rect 38822 280658 58266 280894
rect 58502 280658 58586 280894
rect 58822 280658 78266 280894
rect 78502 280658 78586 280894
rect 78822 280658 98266 280894
rect 98502 280658 98586 280894
rect 98822 280658 118266 280894
rect 118502 280658 118586 280894
rect 118822 280658 138266 280894
rect 138502 280658 138586 280894
rect 138822 280658 158266 280894
rect 158502 280658 158586 280894
rect 158822 280658 178266 280894
rect 178502 280658 178586 280894
rect 178822 280658 198266 280894
rect 198502 280658 198586 280894
rect 198822 280658 218266 280894
rect 218502 280658 218586 280894
rect 218822 280658 238266 280894
rect 238502 280658 238586 280894
rect 238822 280658 258266 280894
rect 258502 280658 258586 280894
rect 258822 280658 278266 280894
rect 278502 280658 278586 280894
rect 278822 280658 298266 280894
rect 298502 280658 298586 280894
rect 298822 280658 318266 280894
rect 318502 280658 318586 280894
rect 318822 280658 338266 280894
rect 338502 280658 338586 280894
rect 338822 280658 358266 280894
rect 358502 280658 358586 280894
rect 358822 280658 378266 280894
rect 378502 280658 378586 280894
rect 378822 280658 398266 280894
rect 398502 280658 398586 280894
rect 398822 280658 418266 280894
rect 418502 280658 418586 280894
rect 418822 280658 438266 280894
rect 438502 280658 438586 280894
rect 438822 280658 458266 280894
rect 458502 280658 458586 280894
rect 458822 280658 478266 280894
rect 478502 280658 478586 280894
rect 478822 280658 498266 280894
rect 498502 280658 498586 280894
rect 498822 280658 518266 280894
rect 518502 280658 518586 280894
rect 518822 280658 538266 280894
rect 538502 280658 538586 280894
rect 538822 280658 558266 280894
rect 558502 280658 558586 280894
rect 558822 280658 578266 280894
rect 578502 280658 578586 280894
rect 578822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 18266 280574
rect 18502 280338 18586 280574
rect 18822 280338 38266 280574
rect 38502 280338 38586 280574
rect 38822 280338 58266 280574
rect 58502 280338 58586 280574
rect 58822 280338 78266 280574
rect 78502 280338 78586 280574
rect 78822 280338 98266 280574
rect 98502 280338 98586 280574
rect 98822 280338 118266 280574
rect 118502 280338 118586 280574
rect 118822 280338 138266 280574
rect 138502 280338 138586 280574
rect 138822 280338 158266 280574
rect 158502 280338 158586 280574
rect 158822 280338 178266 280574
rect 178502 280338 178586 280574
rect 178822 280338 198266 280574
rect 198502 280338 198586 280574
rect 198822 280338 218266 280574
rect 218502 280338 218586 280574
rect 218822 280338 238266 280574
rect 238502 280338 238586 280574
rect 238822 280338 258266 280574
rect 258502 280338 258586 280574
rect 258822 280338 278266 280574
rect 278502 280338 278586 280574
rect 278822 280338 298266 280574
rect 298502 280338 298586 280574
rect 298822 280338 318266 280574
rect 318502 280338 318586 280574
rect 318822 280338 338266 280574
rect 338502 280338 338586 280574
rect 338822 280338 358266 280574
rect 358502 280338 358586 280574
rect 358822 280338 378266 280574
rect 378502 280338 378586 280574
rect 378822 280338 398266 280574
rect 398502 280338 398586 280574
rect 398822 280338 418266 280574
rect 418502 280338 418586 280574
rect 418822 280338 438266 280574
rect 438502 280338 438586 280574
rect 438822 280338 458266 280574
rect 458502 280338 458586 280574
rect 458822 280338 478266 280574
rect 478502 280338 478586 280574
rect 478822 280338 498266 280574
rect 498502 280338 498586 280574
rect 498822 280338 518266 280574
rect 518502 280338 518586 280574
rect 518822 280338 538266 280574
rect 538502 280338 538586 280574
rect 538822 280338 558266 280574
rect 558502 280338 558586 280574
rect 558822 280338 578266 280574
rect 578502 280338 578586 280574
rect 578822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 14546 277174
rect 14782 276938 14866 277174
rect 15102 276938 34546 277174
rect 34782 276938 34866 277174
rect 35102 276938 54546 277174
rect 54782 276938 54866 277174
rect 55102 276938 74546 277174
rect 74782 276938 74866 277174
rect 75102 276938 94546 277174
rect 94782 276938 94866 277174
rect 95102 276938 114546 277174
rect 114782 276938 114866 277174
rect 115102 276938 134546 277174
rect 134782 276938 134866 277174
rect 135102 276938 154546 277174
rect 154782 276938 154866 277174
rect 155102 276938 174546 277174
rect 174782 276938 174866 277174
rect 175102 276938 194546 277174
rect 194782 276938 194866 277174
rect 195102 276938 214546 277174
rect 214782 276938 214866 277174
rect 215102 276938 234546 277174
rect 234782 276938 234866 277174
rect 235102 276938 254546 277174
rect 254782 276938 254866 277174
rect 255102 276938 274546 277174
rect 274782 276938 274866 277174
rect 275102 276938 294546 277174
rect 294782 276938 294866 277174
rect 295102 276938 314546 277174
rect 314782 276938 314866 277174
rect 315102 276938 334546 277174
rect 334782 276938 334866 277174
rect 335102 276938 354546 277174
rect 354782 276938 354866 277174
rect 355102 276938 374546 277174
rect 374782 276938 374866 277174
rect 375102 276938 394546 277174
rect 394782 276938 394866 277174
rect 395102 276938 414546 277174
rect 414782 276938 414866 277174
rect 415102 276938 434546 277174
rect 434782 276938 434866 277174
rect 435102 276938 454546 277174
rect 454782 276938 454866 277174
rect 455102 276938 474546 277174
rect 474782 276938 474866 277174
rect 475102 276938 494546 277174
rect 494782 276938 494866 277174
rect 495102 276938 514546 277174
rect 514782 276938 514866 277174
rect 515102 276938 534546 277174
rect 534782 276938 534866 277174
rect 535102 276938 554546 277174
rect 554782 276938 554866 277174
rect 555102 276938 574546 277174
rect 574782 276938 574866 277174
rect 575102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 14546 276854
rect 14782 276618 14866 276854
rect 15102 276618 34546 276854
rect 34782 276618 34866 276854
rect 35102 276618 54546 276854
rect 54782 276618 54866 276854
rect 55102 276618 74546 276854
rect 74782 276618 74866 276854
rect 75102 276618 94546 276854
rect 94782 276618 94866 276854
rect 95102 276618 114546 276854
rect 114782 276618 114866 276854
rect 115102 276618 134546 276854
rect 134782 276618 134866 276854
rect 135102 276618 154546 276854
rect 154782 276618 154866 276854
rect 155102 276618 174546 276854
rect 174782 276618 174866 276854
rect 175102 276618 194546 276854
rect 194782 276618 194866 276854
rect 195102 276618 214546 276854
rect 214782 276618 214866 276854
rect 215102 276618 234546 276854
rect 234782 276618 234866 276854
rect 235102 276618 254546 276854
rect 254782 276618 254866 276854
rect 255102 276618 274546 276854
rect 274782 276618 274866 276854
rect 275102 276618 294546 276854
rect 294782 276618 294866 276854
rect 295102 276618 314546 276854
rect 314782 276618 314866 276854
rect 315102 276618 334546 276854
rect 334782 276618 334866 276854
rect 335102 276618 354546 276854
rect 354782 276618 354866 276854
rect 355102 276618 374546 276854
rect 374782 276618 374866 276854
rect 375102 276618 394546 276854
rect 394782 276618 394866 276854
rect 395102 276618 414546 276854
rect 414782 276618 414866 276854
rect 415102 276618 434546 276854
rect 434782 276618 434866 276854
rect 435102 276618 454546 276854
rect 454782 276618 454866 276854
rect 455102 276618 474546 276854
rect 474782 276618 474866 276854
rect 475102 276618 494546 276854
rect 494782 276618 494866 276854
rect 495102 276618 514546 276854
rect 514782 276618 514866 276854
rect 515102 276618 534546 276854
rect 534782 276618 534866 276854
rect 535102 276618 554546 276854
rect 554782 276618 554866 276854
rect 555102 276618 574546 276854
rect 574782 276618 574866 276854
rect 575102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 10826 273454
rect 11062 273218 11146 273454
rect 11382 273218 30826 273454
rect 31062 273218 31146 273454
rect 31382 273218 50826 273454
rect 51062 273218 51146 273454
rect 51382 273218 70826 273454
rect 71062 273218 71146 273454
rect 71382 273218 90826 273454
rect 91062 273218 91146 273454
rect 91382 273218 110826 273454
rect 111062 273218 111146 273454
rect 111382 273218 130826 273454
rect 131062 273218 131146 273454
rect 131382 273218 150826 273454
rect 151062 273218 151146 273454
rect 151382 273218 170826 273454
rect 171062 273218 171146 273454
rect 171382 273218 190826 273454
rect 191062 273218 191146 273454
rect 191382 273218 210826 273454
rect 211062 273218 211146 273454
rect 211382 273218 230826 273454
rect 231062 273218 231146 273454
rect 231382 273218 250826 273454
rect 251062 273218 251146 273454
rect 251382 273218 270826 273454
rect 271062 273218 271146 273454
rect 271382 273218 290826 273454
rect 291062 273218 291146 273454
rect 291382 273218 310826 273454
rect 311062 273218 311146 273454
rect 311382 273218 330826 273454
rect 331062 273218 331146 273454
rect 331382 273218 350826 273454
rect 351062 273218 351146 273454
rect 351382 273218 370826 273454
rect 371062 273218 371146 273454
rect 371382 273218 390826 273454
rect 391062 273218 391146 273454
rect 391382 273218 410826 273454
rect 411062 273218 411146 273454
rect 411382 273218 430826 273454
rect 431062 273218 431146 273454
rect 431382 273218 450826 273454
rect 451062 273218 451146 273454
rect 451382 273218 470826 273454
rect 471062 273218 471146 273454
rect 471382 273218 490826 273454
rect 491062 273218 491146 273454
rect 491382 273218 510826 273454
rect 511062 273218 511146 273454
rect 511382 273218 530826 273454
rect 531062 273218 531146 273454
rect 531382 273218 550826 273454
rect 551062 273218 551146 273454
rect 551382 273218 570826 273454
rect 571062 273218 571146 273454
rect 571382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 10826 273134
rect 11062 272898 11146 273134
rect 11382 272898 30826 273134
rect 31062 272898 31146 273134
rect 31382 272898 50826 273134
rect 51062 272898 51146 273134
rect 51382 272898 70826 273134
rect 71062 272898 71146 273134
rect 71382 272898 90826 273134
rect 91062 272898 91146 273134
rect 91382 272898 110826 273134
rect 111062 272898 111146 273134
rect 111382 272898 130826 273134
rect 131062 272898 131146 273134
rect 131382 272898 150826 273134
rect 151062 272898 151146 273134
rect 151382 272898 170826 273134
rect 171062 272898 171146 273134
rect 171382 272898 190826 273134
rect 191062 272898 191146 273134
rect 191382 272898 210826 273134
rect 211062 272898 211146 273134
rect 211382 272898 230826 273134
rect 231062 272898 231146 273134
rect 231382 272898 250826 273134
rect 251062 272898 251146 273134
rect 251382 272898 270826 273134
rect 271062 272898 271146 273134
rect 271382 272898 290826 273134
rect 291062 272898 291146 273134
rect 291382 272898 310826 273134
rect 311062 272898 311146 273134
rect 311382 272898 330826 273134
rect 331062 272898 331146 273134
rect 331382 272898 350826 273134
rect 351062 272898 351146 273134
rect 351382 272898 370826 273134
rect 371062 272898 371146 273134
rect 371382 272898 390826 273134
rect 391062 272898 391146 273134
rect 391382 272898 410826 273134
rect 411062 272898 411146 273134
rect 411382 272898 430826 273134
rect 431062 272898 431146 273134
rect 431382 272898 450826 273134
rect 451062 272898 451146 273134
rect 451382 272898 470826 273134
rect 471062 272898 471146 273134
rect 471382 272898 490826 273134
rect 491062 272898 491146 273134
rect 491382 272898 510826 273134
rect 511062 272898 511146 273134
rect 511382 272898 530826 273134
rect 531062 272898 531146 273134
rect 531382 272898 550826 273134
rect 551062 272898 551146 273134
rect 551382 272898 570826 273134
rect 571062 272898 571146 273134
rect 571382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 11986 266614
rect 12222 266378 12306 266614
rect 12542 266378 31986 266614
rect 32222 266378 32306 266614
rect 32542 266378 51986 266614
rect 52222 266378 52306 266614
rect 52542 266378 71986 266614
rect 72222 266378 72306 266614
rect 72542 266378 91986 266614
rect 92222 266378 92306 266614
rect 92542 266378 111986 266614
rect 112222 266378 112306 266614
rect 112542 266378 131986 266614
rect 132222 266378 132306 266614
rect 132542 266378 151986 266614
rect 152222 266378 152306 266614
rect 152542 266378 171986 266614
rect 172222 266378 172306 266614
rect 172542 266378 191986 266614
rect 192222 266378 192306 266614
rect 192542 266378 211986 266614
rect 212222 266378 212306 266614
rect 212542 266378 231986 266614
rect 232222 266378 232306 266614
rect 232542 266378 251986 266614
rect 252222 266378 252306 266614
rect 252542 266378 271986 266614
rect 272222 266378 272306 266614
rect 272542 266378 291986 266614
rect 292222 266378 292306 266614
rect 292542 266378 311986 266614
rect 312222 266378 312306 266614
rect 312542 266378 331986 266614
rect 332222 266378 332306 266614
rect 332542 266378 351986 266614
rect 352222 266378 352306 266614
rect 352542 266378 371986 266614
rect 372222 266378 372306 266614
rect 372542 266378 391986 266614
rect 392222 266378 392306 266614
rect 392542 266378 411986 266614
rect 412222 266378 412306 266614
rect 412542 266378 431986 266614
rect 432222 266378 432306 266614
rect 432542 266378 451986 266614
rect 452222 266378 452306 266614
rect 452542 266378 471986 266614
rect 472222 266378 472306 266614
rect 472542 266378 491986 266614
rect 492222 266378 492306 266614
rect 492542 266378 511986 266614
rect 512222 266378 512306 266614
rect 512542 266378 531986 266614
rect 532222 266378 532306 266614
rect 532542 266378 551986 266614
rect 552222 266378 552306 266614
rect 552542 266378 571986 266614
rect 572222 266378 572306 266614
rect 572542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 11986 266294
rect 12222 266058 12306 266294
rect 12542 266058 31986 266294
rect 32222 266058 32306 266294
rect 32542 266058 51986 266294
rect 52222 266058 52306 266294
rect 52542 266058 71986 266294
rect 72222 266058 72306 266294
rect 72542 266058 91986 266294
rect 92222 266058 92306 266294
rect 92542 266058 111986 266294
rect 112222 266058 112306 266294
rect 112542 266058 131986 266294
rect 132222 266058 132306 266294
rect 132542 266058 151986 266294
rect 152222 266058 152306 266294
rect 152542 266058 171986 266294
rect 172222 266058 172306 266294
rect 172542 266058 191986 266294
rect 192222 266058 192306 266294
rect 192542 266058 211986 266294
rect 212222 266058 212306 266294
rect 212542 266058 231986 266294
rect 232222 266058 232306 266294
rect 232542 266058 251986 266294
rect 252222 266058 252306 266294
rect 252542 266058 271986 266294
rect 272222 266058 272306 266294
rect 272542 266058 291986 266294
rect 292222 266058 292306 266294
rect 292542 266058 311986 266294
rect 312222 266058 312306 266294
rect 312542 266058 331986 266294
rect 332222 266058 332306 266294
rect 332542 266058 351986 266294
rect 352222 266058 352306 266294
rect 352542 266058 371986 266294
rect 372222 266058 372306 266294
rect 372542 266058 391986 266294
rect 392222 266058 392306 266294
rect 392542 266058 411986 266294
rect 412222 266058 412306 266294
rect 412542 266058 431986 266294
rect 432222 266058 432306 266294
rect 432542 266058 451986 266294
rect 452222 266058 452306 266294
rect 452542 266058 471986 266294
rect 472222 266058 472306 266294
rect 472542 266058 491986 266294
rect 492222 266058 492306 266294
rect 492542 266058 511986 266294
rect 512222 266058 512306 266294
rect 512542 266058 531986 266294
rect 532222 266058 532306 266294
rect 532542 266058 551986 266294
rect 552222 266058 552306 266294
rect 552542 266058 571986 266294
rect 572222 266058 572306 266294
rect 572542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 8266 262894
rect 8502 262658 8586 262894
rect 8822 262658 28266 262894
rect 28502 262658 28586 262894
rect 28822 262658 48266 262894
rect 48502 262658 48586 262894
rect 48822 262658 68266 262894
rect 68502 262658 68586 262894
rect 68822 262658 88266 262894
rect 88502 262658 88586 262894
rect 88822 262658 108266 262894
rect 108502 262658 108586 262894
rect 108822 262658 128266 262894
rect 128502 262658 128586 262894
rect 128822 262658 148266 262894
rect 148502 262658 148586 262894
rect 148822 262658 168266 262894
rect 168502 262658 168586 262894
rect 168822 262658 188266 262894
rect 188502 262658 188586 262894
rect 188822 262658 208266 262894
rect 208502 262658 208586 262894
rect 208822 262658 228266 262894
rect 228502 262658 228586 262894
rect 228822 262658 248266 262894
rect 248502 262658 248586 262894
rect 248822 262658 268266 262894
rect 268502 262658 268586 262894
rect 268822 262658 288266 262894
rect 288502 262658 288586 262894
rect 288822 262658 308266 262894
rect 308502 262658 308586 262894
rect 308822 262658 328266 262894
rect 328502 262658 328586 262894
rect 328822 262658 348266 262894
rect 348502 262658 348586 262894
rect 348822 262658 368266 262894
rect 368502 262658 368586 262894
rect 368822 262658 388266 262894
rect 388502 262658 388586 262894
rect 388822 262658 408266 262894
rect 408502 262658 408586 262894
rect 408822 262658 428266 262894
rect 428502 262658 428586 262894
rect 428822 262658 448266 262894
rect 448502 262658 448586 262894
rect 448822 262658 468266 262894
rect 468502 262658 468586 262894
rect 468822 262658 488266 262894
rect 488502 262658 488586 262894
rect 488822 262658 508266 262894
rect 508502 262658 508586 262894
rect 508822 262658 528266 262894
rect 528502 262658 528586 262894
rect 528822 262658 548266 262894
rect 548502 262658 548586 262894
rect 548822 262658 568266 262894
rect 568502 262658 568586 262894
rect 568822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 8266 262574
rect 8502 262338 8586 262574
rect 8822 262338 28266 262574
rect 28502 262338 28586 262574
rect 28822 262338 48266 262574
rect 48502 262338 48586 262574
rect 48822 262338 68266 262574
rect 68502 262338 68586 262574
rect 68822 262338 88266 262574
rect 88502 262338 88586 262574
rect 88822 262338 108266 262574
rect 108502 262338 108586 262574
rect 108822 262338 128266 262574
rect 128502 262338 128586 262574
rect 128822 262338 148266 262574
rect 148502 262338 148586 262574
rect 148822 262338 168266 262574
rect 168502 262338 168586 262574
rect 168822 262338 188266 262574
rect 188502 262338 188586 262574
rect 188822 262338 208266 262574
rect 208502 262338 208586 262574
rect 208822 262338 228266 262574
rect 228502 262338 228586 262574
rect 228822 262338 248266 262574
rect 248502 262338 248586 262574
rect 248822 262338 268266 262574
rect 268502 262338 268586 262574
rect 268822 262338 288266 262574
rect 288502 262338 288586 262574
rect 288822 262338 308266 262574
rect 308502 262338 308586 262574
rect 308822 262338 328266 262574
rect 328502 262338 328586 262574
rect 328822 262338 348266 262574
rect 348502 262338 348586 262574
rect 348822 262338 368266 262574
rect 368502 262338 368586 262574
rect 368822 262338 388266 262574
rect 388502 262338 388586 262574
rect 388822 262338 408266 262574
rect 408502 262338 408586 262574
rect 408822 262338 428266 262574
rect 428502 262338 428586 262574
rect 428822 262338 448266 262574
rect 448502 262338 448586 262574
rect 448822 262338 468266 262574
rect 468502 262338 468586 262574
rect 468822 262338 488266 262574
rect 488502 262338 488586 262574
rect 488822 262338 508266 262574
rect 508502 262338 508586 262574
rect 508822 262338 528266 262574
rect 528502 262338 528586 262574
rect 528822 262338 548266 262574
rect 548502 262338 548586 262574
rect 548822 262338 568266 262574
rect 568502 262338 568586 262574
rect 568822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 4546 259174
rect 4782 258938 4866 259174
rect 5102 258938 24546 259174
rect 24782 258938 24866 259174
rect 25102 258938 44546 259174
rect 44782 258938 44866 259174
rect 45102 258938 64546 259174
rect 64782 258938 64866 259174
rect 65102 258938 84546 259174
rect 84782 258938 84866 259174
rect 85102 258938 104546 259174
rect 104782 258938 104866 259174
rect 105102 258938 124546 259174
rect 124782 258938 124866 259174
rect 125102 258938 144546 259174
rect 144782 258938 144866 259174
rect 145102 258938 164546 259174
rect 164782 258938 164866 259174
rect 165102 258938 184546 259174
rect 184782 258938 184866 259174
rect 185102 258938 204546 259174
rect 204782 258938 204866 259174
rect 205102 258938 224546 259174
rect 224782 258938 224866 259174
rect 225102 258938 244546 259174
rect 244782 258938 244866 259174
rect 245102 258938 264546 259174
rect 264782 258938 264866 259174
rect 265102 258938 284546 259174
rect 284782 258938 284866 259174
rect 285102 258938 304546 259174
rect 304782 258938 304866 259174
rect 305102 258938 324546 259174
rect 324782 258938 324866 259174
rect 325102 258938 344546 259174
rect 344782 258938 344866 259174
rect 345102 258938 364546 259174
rect 364782 258938 364866 259174
rect 365102 258938 384546 259174
rect 384782 258938 384866 259174
rect 385102 258938 404546 259174
rect 404782 258938 404866 259174
rect 405102 258938 424546 259174
rect 424782 258938 424866 259174
rect 425102 258938 444546 259174
rect 444782 258938 444866 259174
rect 445102 258938 464546 259174
rect 464782 258938 464866 259174
rect 465102 258938 484546 259174
rect 484782 258938 484866 259174
rect 485102 258938 504546 259174
rect 504782 258938 504866 259174
rect 505102 258938 524546 259174
rect 524782 258938 524866 259174
rect 525102 258938 544546 259174
rect 544782 258938 544866 259174
rect 545102 258938 564546 259174
rect 564782 258938 564866 259174
rect 565102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 4546 258854
rect 4782 258618 4866 258854
rect 5102 258618 24546 258854
rect 24782 258618 24866 258854
rect 25102 258618 44546 258854
rect 44782 258618 44866 258854
rect 45102 258618 64546 258854
rect 64782 258618 64866 258854
rect 65102 258618 84546 258854
rect 84782 258618 84866 258854
rect 85102 258618 104546 258854
rect 104782 258618 104866 258854
rect 105102 258618 124546 258854
rect 124782 258618 124866 258854
rect 125102 258618 144546 258854
rect 144782 258618 144866 258854
rect 145102 258618 164546 258854
rect 164782 258618 164866 258854
rect 165102 258618 184546 258854
rect 184782 258618 184866 258854
rect 185102 258618 204546 258854
rect 204782 258618 204866 258854
rect 205102 258618 224546 258854
rect 224782 258618 224866 258854
rect 225102 258618 244546 258854
rect 244782 258618 244866 258854
rect 245102 258618 264546 258854
rect 264782 258618 264866 258854
rect 265102 258618 284546 258854
rect 284782 258618 284866 258854
rect 285102 258618 304546 258854
rect 304782 258618 304866 258854
rect 305102 258618 324546 258854
rect 324782 258618 324866 258854
rect 325102 258618 344546 258854
rect 344782 258618 344866 258854
rect 345102 258618 364546 258854
rect 364782 258618 364866 258854
rect 365102 258618 384546 258854
rect 384782 258618 384866 258854
rect 385102 258618 404546 258854
rect 404782 258618 404866 258854
rect 405102 258618 424546 258854
rect 424782 258618 424866 258854
rect 425102 258618 444546 258854
rect 444782 258618 444866 258854
rect 445102 258618 464546 258854
rect 464782 258618 464866 258854
rect 465102 258618 484546 258854
rect 484782 258618 484866 258854
rect 485102 258618 504546 258854
rect 504782 258618 504866 258854
rect 505102 258618 524546 258854
rect 524782 258618 524866 258854
rect 525102 258618 544546 258854
rect 544782 258618 544866 258854
rect 545102 258618 564546 258854
rect 564782 258618 564866 258854
rect 565102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 826 255454
rect 1062 255218 1146 255454
rect 1382 255218 20826 255454
rect 21062 255218 21146 255454
rect 21382 255218 40826 255454
rect 41062 255218 41146 255454
rect 41382 255218 60826 255454
rect 61062 255218 61146 255454
rect 61382 255218 80826 255454
rect 81062 255218 81146 255454
rect 81382 255218 100826 255454
rect 101062 255218 101146 255454
rect 101382 255218 120826 255454
rect 121062 255218 121146 255454
rect 121382 255218 140826 255454
rect 141062 255218 141146 255454
rect 141382 255218 160826 255454
rect 161062 255218 161146 255454
rect 161382 255218 180826 255454
rect 181062 255218 181146 255454
rect 181382 255218 200826 255454
rect 201062 255218 201146 255454
rect 201382 255218 220826 255454
rect 221062 255218 221146 255454
rect 221382 255218 240826 255454
rect 241062 255218 241146 255454
rect 241382 255218 260826 255454
rect 261062 255218 261146 255454
rect 261382 255218 280826 255454
rect 281062 255218 281146 255454
rect 281382 255218 300826 255454
rect 301062 255218 301146 255454
rect 301382 255218 320826 255454
rect 321062 255218 321146 255454
rect 321382 255218 340826 255454
rect 341062 255218 341146 255454
rect 341382 255218 360826 255454
rect 361062 255218 361146 255454
rect 361382 255218 380826 255454
rect 381062 255218 381146 255454
rect 381382 255218 400826 255454
rect 401062 255218 401146 255454
rect 401382 255218 420826 255454
rect 421062 255218 421146 255454
rect 421382 255218 440826 255454
rect 441062 255218 441146 255454
rect 441382 255218 460826 255454
rect 461062 255218 461146 255454
rect 461382 255218 480826 255454
rect 481062 255218 481146 255454
rect 481382 255218 500826 255454
rect 501062 255218 501146 255454
rect 501382 255218 520826 255454
rect 521062 255218 521146 255454
rect 521382 255218 540826 255454
rect 541062 255218 541146 255454
rect 541382 255218 560826 255454
rect 561062 255218 561146 255454
rect 561382 255218 580826 255454
rect 581062 255218 581146 255454
rect 581382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 826 255134
rect 1062 254898 1146 255134
rect 1382 254898 20826 255134
rect 21062 254898 21146 255134
rect 21382 254898 40826 255134
rect 41062 254898 41146 255134
rect 41382 254898 60826 255134
rect 61062 254898 61146 255134
rect 61382 254898 80826 255134
rect 81062 254898 81146 255134
rect 81382 254898 100826 255134
rect 101062 254898 101146 255134
rect 101382 254898 120826 255134
rect 121062 254898 121146 255134
rect 121382 254898 140826 255134
rect 141062 254898 141146 255134
rect 141382 254898 160826 255134
rect 161062 254898 161146 255134
rect 161382 254898 180826 255134
rect 181062 254898 181146 255134
rect 181382 254898 200826 255134
rect 201062 254898 201146 255134
rect 201382 254898 220826 255134
rect 221062 254898 221146 255134
rect 221382 254898 240826 255134
rect 241062 254898 241146 255134
rect 241382 254898 260826 255134
rect 261062 254898 261146 255134
rect 261382 254898 280826 255134
rect 281062 254898 281146 255134
rect 281382 254898 300826 255134
rect 301062 254898 301146 255134
rect 301382 254898 320826 255134
rect 321062 254898 321146 255134
rect 321382 254898 340826 255134
rect 341062 254898 341146 255134
rect 341382 254898 360826 255134
rect 361062 254898 361146 255134
rect 361382 254898 380826 255134
rect 381062 254898 381146 255134
rect 381382 254898 400826 255134
rect 401062 254898 401146 255134
rect 401382 254898 420826 255134
rect 421062 254898 421146 255134
rect 421382 254898 440826 255134
rect 441062 254898 441146 255134
rect 441382 254898 460826 255134
rect 461062 254898 461146 255134
rect 461382 254898 480826 255134
rect 481062 254898 481146 255134
rect 481382 254898 500826 255134
rect 501062 254898 501146 255134
rect 501382 254898 520826 255134
rect 521062 254898 521146 255134
rect 521382 254898 540826 255134
rect 541062 254898 541146 255134
rect 541382 254898 560826 255134
rect 561062 254898 561146 255134
rect 561382 254898 580826 255134
rect 581062 254898 581146 255134
rect 581382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 21986 248614
rect 22222 248378 22306 248614
rect 22542 248378 41986 248614
rect 42222 248378 42306 248614
rect 42542 248378 61986 248614
rect 62222 248378 62306 248614
rect 62542 248378 81986 248614
rect 82222 248378 82306 248614
rect 82542 248378 101986 248614
rect 102222 248378 102306 248614
rect 102542 248378 121986 248614
rect 122222 248378 122306 248614
rect 122542 248378 141986 248614
rect 142222 248378 142306 248614
rect 142542 248378 161986 248614
rect 162222 248378 162306 248614
rect 162542 248378 181986 248614
rect 182222 248378 182306 248614
rect 182542 248378 201986 248614
rect 202222 248378 202306 248614
rect 202542 248378 221986 248614
rect 222222 248378 222306 248614
rect 222542 248378 241986 248614
rect 242222 248378 242306 248614
rect 242542 248378 261986 248614
rect 262222 248378 262306 248614
rect 262542 248378 281986 248614
rect 282222 248378 282306 248614
rect 282542 248378 301986 248614
rect 302222 248378 302306 248614
rect 302542 248378 321986 248614
rect 322222 248378 322306 248614
rect 322542 248378 341986 248614
rect 342222 248378 342306 248614
rect 342542 248378 361986 248614
rect 362222 248378 362306 248614
rect 362542 248378 381986 248614
rect 382222 248378 382306 248614
rect 382542 248378 401986 248614
rect 402222 248378 402306 248614
rect 402542 248378 421986 248614
rect 422222 248378 422306 248614
rect 422542 248378 441986 248614
rect 442222 248378 442306 248614
rect 442542 248378 461986 248614
rect 462222 248378 462306 248614
rect 462542 248378 481986 248614
rect 482222 248378 482306 248614
rect 482542 248378 501986 248614
rect 502222 248378 502306 248614
rect 502542 248378 521986 248614
rect 522222 248378 522306 248614
rect 522542 248378 541986 248614
rect 542222 248378 542306 248614
rect 542542 248378 561986 248614
rect 562222 248378 562306 248614
rect 562542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 21986 248294
rect 22222 248058 22306 248294
rect 22542 248058 41986 248294
rect 42222 248058 42306 248294
rect 42542 248058 61986 248294
rect 62222 248058 62306 248294
rect 62542 248058 81986 248294
rect 82222 248058 82306 248294
rect 82542 248058 101986 248294
rect 102222 248058 102306 248294
rect 102542 248058 121986 248294
rect 122222 248058 122306 248294
rect 122542 248058 141986 248294
rect 142222 248058 142306 248294
rect 142542 248058 161986 248294
rect 162222 248058 162306 248294
rect 162542 248058 181986 248294
rect 182222 248058 182306 248294
rect 182542 248058 201986 248294
rect 202222 248058 202306 248294
rect 202542 248058 221986 248294
rect 222222 248058 222306 248294
rect 222542 248058 241986 248294
rect 242222 248058 242306 248294
rect 242542 248058 261986 248294
rect 262222 248058 262306 248294
rect 262542 248058 281986 248294
rect 282222 248058 282306 248294
rect 282542 248058 301986 248294
rect 302222 248058 302306 248294
rect 302542 248058 321986 248294
rect 322222 248058 322306 248294
rect 322542 248058 341986 248294
rect 342222 248058 342306 248294
rect 342542 248058 361986 248294
rect 362222 248058 362306 248294
rect 362542 248058 381986 248294
rect 382222 248058 382306 248294
rect 382542 248058 401986 248294
rect 402222 248058 402306 248294
rect 402542 248058 421986 248294
rect 422222 248058 422306 248294
rect 422542 248058 441986 248294
rect 442222 248058 442306 248294
rect 442542 248058 461986 248294
rect 462222 248058 462306 248294
rect 462542 248058 481986 248294
rect 482222 248058 482306 248294
rect 482542 248058 501986 248294
rect 502222 248058 502306 248294
rect 502542 248058 521986 248294
rect 522222 248058 522306 248294
rect 522542 248058 541986 248294
rect 542222 248058 542306 248294
rect 542542 248058 561986 248294
rect 562222 248058 562306 248294
rect 562542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 18266 244894
rect 18502 244658 18586 244894
rect 18822 244658 38266 244894
rect 38502 244658 38586 244894
rect 38822 244658 58266 244894
rect 58502 244658 58586 244894
rect 58822 244658 78266 244894
rect 78502 244658 78586 244894
rect 78822 244658 98266 244894
rect 98502 244658 98586 244894
rect 98822 244658 118266 244894
rect 118502 244658 118586 244894
rect 118822 244658 138266 244894
rect 138502 244658 138586 244894
rect 138822 244658 158266 244894
rect 158502 244658 158586 244894
rect 158822 244658 178266 244894
rect 178502 244658 178586 244894
rect 178822 244658 198266 244894
rect 198502 244658 198586 244894
rect 198822 244658 218266 244894
rect 218502 244658 218586 244894
rect 218822 244658 238266 244894
rect 238502 244658 238586 244894
rect 238822 244658 258266 244894
rect 258502 244658 258586 244894
rect 258822 244658 278266 244894
rect 278502 244658 278586 244894
rect 278822 244658 298266 244894
rect 298502 244658 298586 244894
rect 298822 244658 318266 244894
rect 318502 244658 318586 244894
rect 318822 244658 338266 244894
rect 338502 244658 338586 244894
rect 338822 244658 358266 244894
rect 358502 244658 358586 244894
rect 358822 244658 378266 244894
rect 378502 244658 378586 244894
rect 378822 244658 398266 244894
rect 398502 244658 398586 244894
rect 398822 244658 418266 244894
rect 418502 244658 418586 244894
rect 418822 244658 438266 244894
rect 438502 244658 438586 244894
rect 438822 244658 458266 244894
rect 458502 244658 458586 244894
rect 458822 244658 478266 244894
rect 478502 244658 478586 244894
rect 478822 244658 498266 244894
rect 498502 244658 498586 244894
rect 498822 244658 518266 244894
rect 518502 244658 518586 244894
rect 518822 244658 538266 244894
rect 538502 244658 538586 244894
rect 538822 244658 558266 244894
rect 558502 244658 558586 244894
rect 558822 244658 578266 244894
rect 578502 244658 578586 244894
rect 578822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 18266 244574
rect 18502 244338 18586 244574
rect 18822 244338 38266 244574
rect 38502 244338 38586 244574
rect 38822 244338 58266 244574
rect 58502 244338 58586 244574
rect 58822 244338 78266 244574
rect 78502 244338 78586 244574
rect 78822 244338 98266 244574
rect 98502 244338 98586 244574
rect 98822 244338 118266 244574
rect 118502 244338 118586 244574
rect 118822 244338 138266 244574
rect 138502 244338 138586 244574
rect 138822 244338 158266 244574
rect 158502 244338 158586 244574
rect 158822 244338 178266 244574
rect 178502 244338 178586 244574
rect 178822 244338 198266 244574
rect 198502 244338 198586 244574
rect 198822 244338 218266 244574
rect 218502 244338 218586 244574
rect 218822 244338 238266 244574
rect 238502 244338 238586 244574
rect 238822 244338 258266 244574
rect 258502 244338 258586 244574
rect 258822 244338 278266 244574
rect 278502 244338 278586 244574
rect 278822 244338 298266 244574
rect 298502 244338 298586 244574
rect 298822 244338 318266 244574
rect 318502 244338 318586 244574
rect 318822 244338 338266 244574
rect 338502 244338 338586 244574
rect 338822 244338 358266 244574
rect 358502 244338 358586 244574
rect 358822 244338 378266 244574
rect 378502 244338 378586 244574
rect 378822 244338 398266 244574
rect 398502 244338 398586 244574
rect 398822 244338 418266 244574
rect 418502 244338 418586 244574
rect 418822 244338 438266 244574
rect 438502 244338 438586 244574
rect 438822 244338 458266 244574
rect 458502 244338 458586 244574
rect 458822 244338 478266 244574
rect 478502 244338 478586 244574
rect 478822 244338 498266 244574
rect 498502 244338 498586 244574
rect 498822 244338 518266 244574
rect 518502 244338 518586 244574
rect 518822 244338 538266 244574
rect 538502 244338 538586 244574
rect 538822 244338 558266 244574
rect 558502 244338 558586 244574
rect 558822 244338 578266 244574
rect 578502 244338 578586 244574
rect 578822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 14546 241174
rect 14782 240938 14866 241174
rect 15102 240938 34546 241174
rect 34782 240938 34866 241174
rect 35102 240938 54546 241174
rect 54782 240938 54866 241174
rect 55102 240938 74546 241174
rect 74782 240938 74866 241174
rect 75102 240938 94546 241174
rect 94782 240938 94866 241174
rect 95102 240938 114546 241174
rect 114782 240938 114866 241174
rect 115102 240938 134546 241174
rect 134782 240938 134866 241174
rect 135102 240938 154546 241174
rect 154782 240938 154866 241174
rect 155102 240938 174546 241174
rect 174782 240938 174866 241174
rect 175102 240938 194546 241174
rect 194782 240938 194866 241174
rect 195102 240938 214546 241174
rect 214782 240938 214866 241174
rect 215102 240938 234546 241174
rect 234782 240938 234866 241174
rect 235102 240938 254546 241174
rect 254782 240938 254866 241174
rect 255102 240938 274546 241174
rect 274782 240938 274866 241174
rect 275102 240938 294546 241174
rect 294782 240938 294866 241174
rect 295102 240938 314546 241174
rect 314782 240938 314866 241174
rect 315102 240938 334546 241174
rect 334782 240938 334866 241174
rect 335102 240938 354546 241174
rect 354782 240938 354866 241174
rect 355102 240938 374546 241174
rect 374782 240938 374866 241174
rect 375102 240938 394546 241174
rect 394782 240938 394866 241174
rect 395102 240938 414546 241174
rect 414782 240938 414866 241174
rect 415102 240938 434546 241174
rect 434782 240938 434866 241174
rect 435102 240938 454546 241174
rect 454782 240938 454866 241174
rect 455102 240938 474546 241174
rect 474782 240938 474866 241174
rect 475102 240938 494546 241174
rect 494782 240938 494866 241174
rect 495102 240938 514546 241174
rect 514782 240938 514866 241174
rect 515102 240938 534546 241174
rect 534782 240938 534866 241174
rect 535102 240938 554546 241174
rect 554782 240938 554866 241174
rect 555102 240938 574546 241174
rect 574782 240938 574866 241174
rect 575102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 14546 240854
rect 14782 240618 14866 240854
rect 15102 240618 34546 240854
rect 34782 240618 34866 240854
rect 35102 240618 54546 240854
rect 54782 240618 54866 240854
rect 55102 240618 74546 240854
rect 74782 240618 74866 240854
rect 75102 240618 94546 240854
rect 94782 240618 94866 240854
rect 95102 240618 114546 240854
rect 114782 240618 114866 240854
rect 115102 240618 134546 240854
rect 134782 240618 134866 240854
rect 135102 240618 154546 240854
rect 154782 240618 154866 240854
rect 155102 240618 174546 240854
rect 174782 240618 174866 240854
rect 175102 240618 194546 240854
rect 194782 240618 194866 240854
rect 195102 240618 214546 240854
rect 214782 240618 214866 240854
rect 215102 240618 234546 240854
rect 234782 240618 234866 240854
rect 235102 240618 254546 240854
rect 254782 240618 254866 240854
rect 255102 240618 274546 240854
rect 274782 240618 274866 240854
rect 275102 240618 294546 240854
rect 294782 240618 294866 240854
rect 295102 240618 314546 240854
rect 314782 240618 314866 240854
rect 315102 240618 334546 240854
rect 334782 240618 334866 240854
rect 335102 240618 354546 240854
rect 354782 240618 354866 240854
rect 355102 240618 374546 240854
rect 374782 240618 374866 240854
rect 375102 240618 394546 240854
rect 394782 240618 394866 240854
rect 395102 240618 414546 240854
rect 414782 240618 414866 240854
rect 415102 240618 434546 240854
rect 434782 240618 434866 240854
rect 435102 240618 454546 240854
rect 454782 240618 454866 240854
rect 455102 240618 474546 240854
rect 474782 240618 474866 240854
rect 475102 240618 494546 240854
rect 494782 240618 494866 240854
rect 495102 240618 514546 240854
rect 514782 240618 514866 240854
rect 515102 240618 534546 240854
rect 534782 240618 534866 240854
rect 535102 240618 554546 240854
rect 554782 240618 554866 240854
rect 555102 240618 574546 240854
rect 574782 240618 574866 240854
rect 575102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 10826 237454
rect 11062 237218 11146 237454
rect 11382 237218 30826 237454
rect 31062 237218 31146 237454
rect 31382 237218 50826 237454
rect 51062 237218 51146 237454
rect 51382 237218 70826 237454
rect 71062 237218 71146 237454
rect 71382 237218 90826 237454
rect 91062 237218 91146 237454
rect 91382 237218 110826 237454
rect 111062 237218 111146 237454
rect 111382 237218 130826 237454
rect 131062 237218 131146 237454
rect 131382 237218 150826 237454
rect 151062 237218 151146 237454
rect 151382 237218 170826 237454
rect 171062 237218 171146 237454
rect 171382 237218 190826 237454
rect 191062 237218 191146 237454
rect 191382 237218 210826 237454
rect 211062 237218 211146 237454
rect 211382 237218 230826 237454
rect 231062 237218 231146 237454
rect 231382 237218 250826 237454
rect 251062 237218 251146 237454
rect 251382 237218 270826 237454
rect 271062 237218 271146 237454
rect 271382 237218 290826 237454
rect 291062 237218 291146 237454
rect 291382 237218 310826 237454
rect 311062 237218 311146 237454
rect 311382 237218 330826 237454
rect 331062 237218 331146 237454
rect 331382 237218 350826 237454
rect 351062 237218 351146 237454
rect 351382 237218 370826 237454
rect 371062 237218 371146 237454
rect 371382 237218 390826 237454
rect 391062 237218 391146 237454
rect 391382 237218 410826 237454
rect 411062 237218 411146 237454
rect 411382 237218 430826 237454
rect 431062 237218 431146 237454
rect 431382 237218 450826 237454
rect 451062 237218 451146 237454
rect 451382 237218 470826 237454
rect 471062 237218 471146 237454
rect 471382 237218 490826 237454
rect 491062 237218 491146 237454
rect 491382 237218 510826 237454
rect 511062 237218 511146 237454
rect 511382 237218 530826 237454
rect 531062 237218 531146 237454
rect 531382 237218 550826 237454
rect 551062 237218 551146 237454
rect 551382 237218 570826 237454
rect 571062 237218 571146 237454
rect 571382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 10826 237134
rect 11062 236898 11146 237134
rect 11382 236898 30826 237134
rect 31062 236898 31146 237134
rect 31382 236898 50826 237134
rect 51062 236898 51146 237134
rect 51382 236898 70826 237134
rect 71062 236898 71146 237134
rect 71382 236898 90826 237134
rect 91062 236898 91146 237134
rect 91382 236898 110826 237134
rect 111062 236898 111146 237134
rect 111382 236898 130826 237134
rect 131062 236898 131146 237134
rect 131382 236898 150826 237134
rect 151062 236898 151146 237134
rect 151382 236898 170826 237134
rect 171062 236898 171146 237134
rect 171382 236898 190826 237134
rect 191062 236898 191146 237134
rect 191382 236898 210826 237134
rect 211062 236898 211146 237134
rect 211382 236898 230826 237134
rect 231062 236898 231146 237134
rect 231382 236898 250826 237134
rect 251062 236898 251146 237134
rect 251382 236898 270826 237134
rect 271062 236898 271146 237134
rect 271382 236898 290826 237134
rect 291062 236898 291146 237134
rect 291382 236898 310826 237134
rect 311062 236898 311146 237134
rect 311382 236898 330826 237134
rect 331062 236898 331146 237134
rect 331382 236898 350826 237134
rect 351062 236898 351146 237134
rect 351382 236898 370826 237134
rect 371062 236898 371146 237134
rect 371382 236898 390826 237134
rect 391062 236898 391146 237134
rect 391382 236898 410826 237134
rect 411062 236898 411146 237134
rect 411382 236898 430826 237134
rect 431062 236898 431146 237134
rect 431382 236898 450826 237134
rect 451062 236898 451146 237134
rect 451382 236898 470826 237134
rect 471062 236898 471146 237134
rect 471382 236898 490826 237134
rect 491062 236898 491146 237134
rect 491382 236898 510826 237134
rect 511062 236898 511146 237134
rect 511382 236898 530826 237134
rect 531062 236898 531146 237134
rect 531382 236898 550826 237134
rect 551062 236898 551146 237134
rect 551382 236898 570826 237134
rect 571062 236898 571146 237134
rect 571382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 11986 230614
rect 12222 230378 12306 230614
rect 12542 230378 31986 230614
rect 32222 230378 32306 230614
rect 32542 230378 51986 230614
rect 52222 230378 52306 230614
rect 52542 230378 71986 230614
rect 72222 230378 72306 230614
rect 72542 230378 91986 230614
rect 92222 230378 92306 230614
rect 92542 230378 111986 230614
rect 112222 230378 112306 230614
rect 112542 230378 131986 230614
rect 132222 230378 132306 230614
rect 132542 230378 151986 230614
rect 152222 230378 152306 230614
rect 152542 230378 171986 230614
rect 172222 230378 172306 230614
rect 172542 230378 191986 230614
rect 192222 230378 192306 230614
rect 192542 230378 211986 230614
rect 212222 230378 212306 230614
rect 212542 230378 231986 230614
rect 232222 230378 232306 230614
rect 232542 230378 251986 230614
rect 252222 230378 252306 230614
rect 252542 230378 271986 230614
rect 272222 230378 272306 230614
rect 272542 230378 291986 230614
rect 292222 230378 292306 230614
rect 292542 230378 311986 230614
rect 312222 230378 312306 230614
rect 312542 230378 331986 230614
rect 332222 230378 332306 230614
rect 332542 230378 351986 230614
rect 352222 230378 352306 230614
rect 352542 230378 371986 230614
rect 372222 230378 372306 230614
rect 372542 230378 391986 230614
rect 392222 230378 392306 230614
rect 392542 230378 411986 230614
rect 412222 230378 412306 230614
rect 412542 230378 431986 230614
rect 432222 230378 432306 230614
rect 432542 230378 451986 230614
rect 452222 230378 452306 230614
rect 452542 230378 471986 230614
rect 472222 230378 472306 230614
rect 472542 230378 491986 230614
rect 492222 230378 492306 230614
rect 492542 230378 511986 230614
rect 512222 230378 512306 230614
rect 512542 230378 531986 230614
rect 532222 230378 532306 230614
rect 532542 230378 551986 230614
rect 552222 230378 552306 230614
rect 552542 230378 571986 230614
rect 572222 230378 572306 230614
rect 572542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 11986 230294
rect 12222 230058 12306 230294
rect 12542 230058 31986 230294
rect 32222 230058 32306 230294
rect 32542 230058 51986 230294
rect 52222 230058 52306 230294
rect 52542 230058 71986 230294
rect 72222 230058 72306 230294
rect 72542 230058 91986 230294
rect 92222 230058 92306 230294
rect 92542 230058 111986 230294
rect 112222 230058 112306 230294
rect 112542 230058 131986 230294
rect 132222 230058 132306 230294
rect 132542 230058 151986 230294
rect 152222 230058 152306 230294
rect 152542 230058 171986 230294
rect 172222 230058 172306 230294
rect 172542 230058 191986 230294
rect 192222 230058 192306 230294
rect 192542 230058 211986 230294
rect 212222 230058 212306 230294
rect 212542 230058 231986 230294
rect 232222 230058 232306 230294
rect 232542 230058 251986 230294
rect 252222 230058 252306 230294
rect 252542 230058 271986 230294
rect 272222 230058 272306 230294
rect 272542 230058 291986 230294
rect 292222 230058 292306 230294
rect 292542 230058 311986 230294
rect 312222 230058 312306 230294
rect 312542 230058 331986 230294
rect 332222 230058 332306 230294
rect 332542 230058 351986 230294
rect 352222 230058 352306 230294
rect 352542 230058 371986 230294
rect 372222 230058 372306 230294
rect 372542 230058 391986 230294
rect 392222 230058 392306 230294
rect 392542 230058 411986 230294
rect 412222 230058 412306 230294
rect 412542 230058 431986 230294
rect 432222 230058 432306 230294
rect 432542 230058 451986 230294
rect 452222 230058 452306 230294
rect 452542 230058 471986 230294
rect 472222 230058 472306 230294
rect 472542 230058 491986 230294
rect 492222 230058 492306 230294
rect 492542 230058 511986 230294
rect 512222 230058 512306 230294
rect 512542 230058 531986 230294
rect 532222 230058 532306 230294
rect 532542 230058 551986 230294
rect 552222 230058 552306 230294
rect 552542 230058 571986 230294
rect 572222 230058 572306 230294
rect 572542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 8266 226894
rect 8502 226658 8586 226894
rect 8822 226658 28266 226894
rect 28502 226658 28586 226894
rect 28822 226658 48266 226894
rect 48502 226658 48586 226894
rect 48822 226658 68266 226894
rect 68502 226658 68586 226894
rect 68822 226658 88266 226894
rect 88502 226658 88586 226894
rect 88822 226658 108266 226894
rect 108502 226658 108586 226894
rect 108822 226658 128266 226894
rect 128502 226658 128586 226894
rect 128822 226658 148266 226894
rect 148502 226658 148586 226894
rect 148822 226658 168266 226894
rect 168502 226658 168586 226894
rect 168822 226658 188266 226894
rect 188502 226658 188586 226894
rect 188822 226658 208266 226894
rect 208502 226658 208586 226894
rect 208822 226658 228266 226894
rect 228502 226658 228586 226894
rect 228822 226658 248266 226894
rect 248502 226658 248586 226894
rect 248822 226658 268266 226894
rect 268502 226658 268586 226894
rect 268822 226658 288266 226894
rect 288502 226658 288586 226894
rect 288822 226658 308266 226894
rect 308502 226658 308586 226894
rect 308822 226658 328266 226894
rect 328502 226658 328586 226894
rect 328822 226658 348266 226894
rect 348502 226658 348586 226894
rect 348822 226658 368266 226894
rect 368502 226658 368586 226894
rect 368822 226658 388266 226894
rect 388502 226658 388586 226894
rect 388822 226658 408266 226894
rect 408502 226658 408586 226894
rect 408822 226658 428266 226894
rect 428502 226658 428586 226894
rect 428822 226658 448266 226894
rect 448502 226658 448586 226894
rect 448822 226658 468266 226894
rect 468502 226658 468586 226894
rect 468822 226658 488266 226894
rect 488502 226658 488586 226894
rect 488822 226658 508266 226894
rect 508502 226658 508586 226894
rect 508822 226658 528266 226894
rect 528502 226658 528586 226894
rect 528822 226658 548266 226894
rect 548502 226658 548586 226894
rect 548822 226658 568266 226894
rect 568502 226658 568586 226894
rect 568822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 8266 226574
rect 8502 226338 8586 226574
rect 8822 226338 28266 226574
rect 28502 226338 28586 226574
rect 28822 226338 48266 226574
rect 48502 226338 48586 226574
rect 48822 226338 68266 226574
rect 68502 226338 68586 226574
rect 68822 226338 88266 226574
rect 88502 226338 88586 226574
rect 88822 226338 108266 226574
rect 108502 226338 108586 226574
rect 108822 226338 128266 226574
rect 128502 226338 128586 226574
rect 128822 226338 148266 226574
rect 148502 226338 148586 226574
rect 148822 226338 168266 226574
rect 168502 226338 168586 226574
rect 168822 226338 188266 226574
rect 188502 226338 188586 226574
rect 188822 226338 208266 226574
rect 208502 226338 208586 226574
rect 208822 226338 228266 226574
rect 228502 226338 228586 226574
rect 228822 226338 248266 226574
rect 248502 226338 248586 226574
rect 248822 226338 268266 226574
rect 268502 226338 268586 226574
rect 268822 226338 288266 226574
rect 288502 226338 288586 226574
rect 288822 226338 308266 226574
rect 308502 226338 308586 226574
rect 308822 226338 328266 226574
rect 328502 226338 328586 226574
rect 328822 226338 348266 226574
rect 348502 226338 348586 226574
rect 348822 226338 368266 226574
rect 368502 226338 368586 226574
rect 368822 226338 388266 226574
rect 388502 226338 388586 226574
rect 388822 226338 408266 226574
rect 408502 226338 408586 226574
rect 408822 226338 428266 226574
rect 428502 226338 428586 226574
rect 428822 226338 448266 226574
rect 448502 226338 448586 226574
rect 448822 226338 468266 226574
rect 468502 226338 468586 226574
rect 468822 226338 488266 226574
rect 488502 226338 488586 226574
rect 488822 226338 508266 226574
rect 508502 226338 508586 226574
rect 508822 226338 528266 226574
rect 528502 226338 528586 226574
rect 528822 226338 548266 226574
rect 548502 226338 548586 226574
rect 548822 226338 568266 226574
rect 568502 226338 568586 226574
rect 568822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 4546 223174
rect 4782 222938 4866 223174
rect 5102 222938 24546 223174
rect 24782 222938 24866 223174
rect 25102 222938 44546 223174
rect 44782 222938 44866 223174
rect 45102 222938 64546 223174
rect 64782 222938 64866 223174
rect 65102 222938 84546 223174
rect 84782 222938 84866 223174
rect 85102 222938 104546 223174
rect 104782 222938 104866 223174
rect 105102 222938 124546 223174
rect 124782 222938 124866 223174
rect 125102 222938 144546 223174
rect 144782 222938 144866 223174
rect 145102 222938 164546 223174
rect 164782 222938 164866 223174
rect 165102 222938 184546 223174
rect 184782 222938 184866 223174
rect 185102 222938 204546 223174
rect 204782 222938 204866 223174
rect 205102 222938 224546 223174
rect 224782 222938 224866 223174
rect 225102 222938 244546 223174
rect 244782 222938 244866 223174
rect 245102 222938 264546 223174
rect 264782 222938 264866 223174
rect 265102 222938 284546 223174
rect 284782 222938 284866 223174
rect 285102 222938 304546 223174
rect 304782 222938 304866 223174
rect 305102 222938 324546 223174
rect 324782 222938 324866 223174
rect 325102 222938 344546 223174
rect 344782 222938 344866 223174
rect 345102 222938 364546 223174
rect 364782 222938 364866 223174
rect 365102 222938 384546 223174
rect 384782 222938 384866 223174
rect 385102 222938 404546 223174
rect 404782 222938 404866 223174
rect 405102 222938 424546 223174
rect 424782 222938 424866 223174
rect 425102 222938 444546 223174
rect 444782 222938 444866 223174
rect 445102 222938 464546 223174
rect 464782 222938 464866 223174
rect 465102 222938 484546 223174
rect 484782 222938 484866 223174
rect 485102 222938 504546 223174
rect 504782 222938 504866 223174
rect 505102 222938 524546 223174
rect 524782 222938 524866 223174
rect 525102 222938 544546 223174
rect 544782 222938 544866 223174
rect 545102 222938 564546 223174
rect 564782 222938 564866 223174
rect 565102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 4546 222854
rect 4782 222618 4866 222854
rect 5102 222618 24546 222854
rect 24782 222618 24866 222854
rect 25102 222618 44546 222854
rect 44782 222618 44866 222854
rect 45102 222618 64546 222854
rect 64782 222618 64866 222854
rect 65102 222618 84546 222854
rect 84782 222618 84866 222854
rect 85102 222618 104546 222854
rect 104782 222618 104866 222854
rect 105102 222618 124546 222854
rect 124782 222618 124866 222854
rect 125102 222618 144546 222854
rect 144782 222618 144866 222854
rect 145102 222618 164546 222854
rect 164782 222618 164866 222854
rect 165102 222618 184546 222854
rect 184782 222618 184866 222854
rect 185102 222618 204546 222854
rect 204782 222618 204866 222854
rect 205102 222618 224546 222854
rect 224782 222618 224866 222854
rect 225102 222618 244546 222854
rect 244782 222618 244866 222854
rect 245102 222618 264546 222854
rect 264782 222618 264866 222854
rect 265102 222618 284546 222854
rect 284782 222618 284866 222854
rect 285102 222618 304546 222854
rect 304782 222618 304866 222854
rect 305102 222618 324546 222854
rect 324782 222618 324866 222854
rect 325102 222618 344546 222854
rect 344782 222618 344866 222854
rect 345102 222618 364546 222854
rect 364782 222618 364866 222854
rect 365102 222618 384546 222854
rect 384782 222618 384866 222854
rect 385102 222618 404546 222854
rect 404782 222618 404866 222854
rect 405102 222618 424546 222854
rect 424782 222618 424866 222854
rect 425102 222618 444546 222854
rect 444782 222618 444866 222854
rect 445102 222618 464546 222854
rect 464782 222618 464866 222854
rect 465102 222618 484546 222854
rect 484782 222618 484866 222854
rect 485102 222618 504546 222854
rect 504782 222618 504866 222854
rect 505102 222618 524546 222854
rect 524782 222618 524866 222854
rect 525102 222618 544546 222854
rect 544782 222618 544866 222854
rect 545102 222618 564546 222854
rect 564782 222618 564866 222854
rect 565102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 826 219454
rect 1062 219218 1146 219454
rect 1382 219218 20826 219454
rect 21062 219218 21146 219454
rect 21382 219218 40826 219454
rect 41062 219218 41146 219454
rect 41382 219218 60826 219454
rect 61062 219218 61146 219454
rect 61382 219218 80826 219454
rect 81062 219218 81146 219454
rect 81382 219218 100826 219454
rect 101062 219218 101146 219454
rect 101382 219218 120826 219454
rect 121062 219218 121146 219454
rect 121382 219218 140826 219454
rect 141062 219218 141146 219454
rect 141382 219218 160826 219454
rect 161062 219218 161146 219454
rect 161382 219218 180826 219454
rect 181062 219218 181146 219454
rect 181382 219218 200826 219454
rect 201062 219218 201146 219454
rect 201382 219218 220826 219454
rect 221062 219218 221146 219454
rect 221382 219218 240826 219454
rect 241062 219218 241146 219454
rect 241382 219218 260826 219454
rect 261062 219218 261146 219454
rect 261382 219218 280826 219454
rect 281062 219218 281146 219454
rect 281382 219218 300826 219454
rect 301062 219218 301146 219454
rect 301382 219218 320826 219454
rect 321062 219218 321146 219454
rect 321382 219218 340826 219454
rect 341062 219218 341146 219454
rect 341382 219218 360826 219454
rect 361062 219218 361146 219454
rect 361382 219218 380826 219454
rect 381062 219218 381146 219454
rect 381382 219218 400826 219454
rect 401062 219218 401146 219454
rect 401382 219218 420826 219454
rect 421062 219218 421146 219454
rect 421382 219218 440826 219454
rect 441062 219218 441146 219454
rect 441382 219218 460826 219454
rect 461062 219218 461146 219454
rect 461382 219218 480826 219454
rect 481062 219218 481146 219454
rect 481382 219218 500826 219454
rect 501062 219218 501146 219454
rect 501382 219218 520826 219454
rect 521062 219218 521146 219454
rect 521382 219218 540826 219454
rect 541062 219218 541146 219454
rect 541382 219218 560826 219454
rect 561062 219218 561146 219454
rect 561382 219218 580826 219454
rect 581062 219218 581146 219454
rect 581382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 826 219134
rect 1062 218898 1146 219134
rect 1382 218898 20826 219134
rect 21062 218898 21146 219134
rect 21382 218898 40826 219134
rect 41062 218898 41146 219134
rect 41382 218898 60826 219134
rect 61062 218898 61146 219134
rect 61382 218898 80826 219134
rect 81062 218898 81146 219134
rect 81382 218898 100826 219134
rect 101062 218898 101146 219134
rect 101382 218898 120826 219134
rect 121062 218898 121146 219134
rect 121382 218898 140826 219134
rect 141062 218898 141146 219134
rect 141382 218898 160826 219134
rect 161062 218898 161146 219134
rect 161382 218898 180826 219134
rect 181062 218898 181146 219134
rect 181382 218898 200826 219134
rect 201062 218898 201146 219134
rect 201382 218898 220826 219134
rect 221062 218898 221146 219134
rect 221382 218898 240826 219134
rect 241062 218898 241146 219134
rect 241382 218898 260826 219134
rect 261062 218898 261146 219134
rect 261382 218898 280826 219134
rect 281062 218898 281146 219134
rect 281382 218898 300826 219134
rect 301062 218898 301146 219134
rect 301382 218898 320826 219134
rect 321062 218898 321146 219134
rect 321382 218898 340826 219134
rect 341062 218898 341146 219134
rect 341382 218898 360826 219134
rect 361062 218898 361146 219134
rect 361382 218898 380826 219134
rect 381062 218898 381146 219134
rect 381382 218898 400826 219134
rect 401062 218898 401146 219134
rect 401382 218898 420826 219134
rect 421062 218898 421146 219134
rect 421382 218898 440826 219134
rect 441062 218898 441146 219134
rect 441382 218898 460826 219134
rect 461062 218898 461146 219134
rect 461382 218898 480826 219134
rect 481062 218898 481146 219134
rect 481382 218898 500826 219134
rect 501062 218898 501146 219134
rect 501382 218898 520826 219134
rect 521062 218898 521146 219134
rect 521382 218898 540826 219134
rect 541062 218898 541146 219134
rect 541382 218898 560826 219134
rect 561062 218898 561146 219134
rect 561382 218898 580826 219134
rect 581062 218898 581146 219134
rect 581382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 21986 212614
rect 22222 212378 22306 212614
rect 22542 212378 41986 212614
rect 42222 212378 42306 212614
rect 42542 212378 61986 212614
rect 62222 212378 62306 212614
rect 62542 212378 81986 212614
rect 82222 212378 82306 212614
rect 82542 212378 101986 212614
rect 102222 212378 102306 212614
rect 102542 212378 121986 212614
rect 122222 212378 122306 212614
rect 122542 212378 141986 212614
rect 142222 212378 142306 212614
rect 142542 212378 161986 212614
rect 162222 212378 162306 212614
rect 162542 212378 181986 212614
rect 182222 212378 182306 212614
rect 182542 212378 201986 212614
rect 202222 212378 202306 212614
rect 202542 212378 221986 212614
rect 222222 212378 222306 212614
rect 222542 212378 241986 212614
rect 242222 212378 242306 212614
rect 242542 212378 261986 212614
rect 262222 212378 262306 212614
rect 262542 212378 281986 212614
rect 282222 212378 282306 212614
rect 282542 212378 301986 212614
rect 302222 212378 302306 212614
rect 302542 212378 321986 212614
rect 322222 212378 322306 212614
rect 322542 212378 341986 212614
rect 342222 212378 342306 212614
rect 342542 212378 361986 212614
rect 362222 212378 362306 212614
rect 362542 212378 381986 212614
rect 382222 212378 382306 212614
rect 382542 212378 401986 212614
rect 402222 212378 402306 212614
rect 402542 212378 421986 212614
rect 422222 212378 422306 212614
rect 422542 212378 441986 212614
rect 442222 212378 442306 212614
rect 442542 212378 461986 212614
rect 462222 212378 462306 212614
rect 462542 212378 481986 212614
rect 482222 212378 482306 212614
rect 482542 212378 501986 212614
rect 502222 212378 502306 212614
rect 502542 212378 521986 212614
rect 522222 212378 522306 212614
rect 522542 212378 541986 212614
rect 542222 212378 542306 212614
rect 542542 212378 561986 212614
rect 562222 212378 562306 212614
rect 562542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 21986 212294
rect 22222 212058 22306 212294
rect 22542 212058 41986 212294
rect 42222 212058 42306 212294
rect 42542 212058 61986 212294
rect 62222 212058 62306 212294
rect 62542 212058 81986 212294
rect 82222 212058 82306 212294
rect 82542 212058 101986 212294
rect 102222 212058 102306 212294
rect 102542 212058 121986 212294
rect 122222 212058 122306 212294
rect 122542 212058 141986 212294
rect 142222 212058 142306 212294
rect 142542 212058 161986 212294
rect 162222 212058 162306 212294
rect 162542 212058 181986 212294
rect 182222 212058 182306 212294
rect 182542 212058 201986 212294
rect 202222 212058 202306 212294
rect 202542 212058 221986 212294
rect 222222 212058 222306 212294
rect 222542 212058 241986 212294
rect 242222 212058 242306 212294
rect 242542 212058 261986 212294
rect 262222 212058 262306 212294
rect 262542 212058 281986 212294
rect 282222 212058 282306 212294
rect 282542 212058 301986 212294
rect 302222 212058 302306 212294
rect 302542 212058 321986 212294
rect 322222 212058 322306 212294
rect 322542 212058 341986 212294
rect 342222 212058 342306 212294
rect 342542 212058 361986 212294
rect 362222 212058 362306 212294
rect 362542 212058 381986 212294
rect 382222 212058 382306 212294
rect 382542 212058 401986 212294
rect 402222 212058 402306 212294
rect 402542 212058 421986 212294
rect 422222 212058 422306 212294
rect 422542 212058 441986 212294
rect 442222 212058 442306 212294
rect 442542 212058 461986 212294
rect 462222 212058 462306 212294
rect 462542 212058 481986 212294
rect 482222 212058 482306 212294
rect 482542 212058 501986 212294
rect 502222 212058 502306 212294
rect 502542 212058 521986 212294
rect 522222 212058 522306 212294
rect 522542 212058 541986 212294
rect 542222 212058 542306 212294
rect 542542 212058 561986 212294
rect 562222 212058 562306 212294
rect 562542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 18266 208894
rect 18502 208658 18586 208894
rect 18822 208658 38266 208894
rect 38502 208658 38586 208894
rect 38822 208658 58266 208894
rect 58502 208658 58586 208894
rect 58822 208658 78266 208894
rect 78502 208658 78586 208894
rect 78822 208658 98266 208894
rect 98502 208658 98586 208894
rect 98822 208658 118266 208894
rect 118502 208658 118586 208894
rect 118822 208658 138266 208894
rect 138502 208658 138586 208894
rect 138822 208658 158266 208894
rect 158502 208658 158586 208894
rect 158822 208658 178266 208894
rect 178502 208658 178586 208894
rect 178822 208658 198266 208894
rect 198502 208658 198586 208894
rect 198822 208658 218266 208894
rect 218502 208658 218586 208894
rect 218822 208658 238266 208894
rect 238502 208658 238586 208894
rect 238822 208658 258266 208894
rect 258502 208658 258586 208894
rect 258822 208658 278266 208894
rect 278502 208658 278586 208894
rect 278822 208658 298266 208894
rect 298502 208658 298586 208894
rect 298822 208658 318266 208894
rect 318502 208658 318586 208894
rect 318822 208658 338266 208894
rect 338502 208658 338586 208894
rect 338822 208658 358266 208894
rect 358502 208658 358586 208894
rect 358822 208658 378266 208894
rect 378502 208658 378586 208894
rect 378822 208658 398266 208894
rect 398502 208658 398586 208894
rect 398822 208658 418266 208894
rect 418502 208658 418586 208894
rect 418822 208658 438266 208894
rect 438502 208658 438586 208894
rect 438822 208658 458266 208894
rect 458502 208658 458586 208894
rect 458822 208658 478266 208894
rect 478502 208658 478586 208894
rect 478822 208658 498266 208894
rect 498502 208658 498586 208894
rect 498822 208658 518266 208894
rect 518502 208658 518586 208894
rect 518822 208658 538266 208894
rect 538502 208658 538586 208894
rect 538822 208658 558266 208894
rect 558502 208658 558586 208894
rect 558822 208658 578266 208894
rect 578502 208658 578586 208894
rect 578822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 18266 208574
rect 18502 208338 18586 208574
rect 18822 208338 38266 208574
rect 38502 208338 38586 208574
rect 38822 208338 58266 208574
rect 58502 208338 58586 208574
rect 58822 208338 78266 208574
rect 78502 208338 78586 208574
rect 78822 208338 98266 208574
rect 98502 208338 98586 208574
rect 98822 208338 118266 208574
rect 118502 208338 118586 208574
rect 118822 208338 138266 208574
rect 138502 208338 138586 208574
rect 138822 208338 158266 208574
rect 158502 208338 158586 208574
rect 158822 208338 178266 208574
rect 178502 208338 178586 208574
rect 178822 208338 198266 208574
rect 198502 208338 198586 208574
rect 198822 208338 218266 208574
rect 218502 208338 218586 208574
rect 218822 208338 238266 208574
rect 238502 208338 238586 208574
rect 238822 208338 258266 208574
rect 258502 208338 258586 208574
rect 258822 208338 278266 208574
rect 278502 208338 278586 208574
rect 278822 208338 298266 208574
rect 298502 208338 298586 208574
rect 298822 208338 318266 208574
rect 318502 208338 318586 208574
rect 318822 208338 338266 208574
rect 338502 208338 338586 208574
rect 338822 208338 358266 208574
rect 358502 208338 358586 208574
rect 358822 208338 378266 208574
rect 378502 208338 378586 208574
rect 378822 208338 398266 208574
rect 398502 208338 398586 208574
rect 398822 208338 418266 208574
rect 418502 208338 418586 208574
rect 418822 208338 438266 208574
rect 438502 208338 438586 208574
rect 438822 208338 458266 208574
rect 458502 208338 458586 208574
rect 458822 208338 478266 208574
rect 478502 208338 478586 208574
rect 478822 208338 498266 208574
rect 498502 208338 498586 208574
rect 498822 208338 518266 208574
rect 518502 208338 518586 208574
rect 518822 208338 538266 208574
rect 538502 208338 538586 208574
rect 538822 208338 558266 208574
rect 558502 208338 558586 208574
rect 558822 208338 578266 208574
rect 578502 208338 578586 208574
rect 578822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 14546 205174
rect 14782 204938 14866 205174
rect 15102 204938 34546 205174
rect 34782 204938 34866 205174
rect 35102 204938 54546 205174
rect 54782 204938 54866 205174
rect 55102 204938 74546 205174
rect 74782 204938 74866 205174
rect 75102 204938 94546 205174
rect 94782 204938 94866 205174
rect 95102 204938 114546 205174
rect 114782 204938 114866 205174
rect 115102 204938 134546 205174
rect 134782 204938 134866 205174
rect 135102 204938 154546 205174
rect 154782 204938 154866 205174
rect 155102 204938 174546 205174
rect 174782 204938 174866 205174
rect 175102 204938 194546 205174
rect 194782 204938 194866 205174
rect 195102 204938 214546 205174
rect 214782 204938 214866 205174
rect 215102 204938 234546 205174
rect 234782 204938 234866 205174
rect 235102 204938 254546 205174
rect 254782 204938 254866 205174
rect 255102 204938 274546 205174
rect 274782 204938 274866 205174
rect 275102 204938 294546 205174
rect 294782 204938 294866 205174
rect 295102 204938 314546 205174
rect 314782 204938 314866 205174
rect 315102 204938 334546 205174
rect 334782 204938 334866 205174
rect 335102 204938 354546 205174
rect 354782 204938 354866 205174
rect 355102 204938 374546 205174
rect 374782 204938 374866 205174
rect 375102 204938 394546 205174
rect 394782 204938 394866 205174
rect 395102 204938 414546 205174
rect 414782 204938 414866 205174
rect 415102 204938 434546 205174
rect 434782 204938 434866 205174
rect 435102 204938 454546 205174
rect 454782 204938 454866 205174
rect 455102 204938 474546 205174
rect 474782 204938 474866 205174
rect 475102 204938 494546 205174
rect 494782 204938 494866 205174
rect 495102 204938 514546 205174
rect 514782 204938 514866 205174
rect 515102 204938 534546 205174
rect 534782 204938 534866 205174
rect 535102 204938 554546 205174
rect 554782 204938 554866 205174
rect 555102 204938 574546 205174
rect 574782 204938 574866 205174
rect 575102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 14546 204854
rect 14782 204618 14866 204854
rect 15102 204618 34546 204854
rect 34782 204618 34866 204854
rect 35102 204618 54546 204854
rect 54782 204618 54866 204854
rect 55102 204618 74546 204854
rect 74782 204618 74866 204854
rect 75102 204618 94546 204854
rect 94782 204618 94866 204854
rect 95102 204618 114546 204854
rect 114782 204618 114866 204854
rect 115102 204618 134546 204854
rect 134782 204618 134866 204854
rect 135102 204618 154546 204854
rect 154782 204618 154866 204854
rect 155102 204618 174546 204854
rect 174782 204618 174866 204854
rect 175102 204618 194546 204854
rect 194782 204618 194866 204854
rect 195102 204618 214546 204854
rect 214782 204618 214866 204854
rect 215102 204618 234546 204854
rect 234782 204618 234866 204854
rect 235102 204618 254546 204854
rect 254782 204618 254866 204854
rect 255102 204618 274546 204854
rect 274782 204618 274866 204854
rect 275102 204618 294546 204854
rect 294782 204618 294866 204854
rect 295102 204618 314546 204854
rect 314782 204618 314866 204854
rect 315102 204618 334546 204854
rect 334782 204618 334866 204854
rect 335102 204618 354546 204854
rect 354782 204618 354866 204854
rect 355102 204618 374546 204854
rect 374782 204618 374866 204854
rect 375102 204618 394546 204854
rect 394782 204618 394866 204854
rect 395102 204618 414546 204854
rect 414782 204618 414866 204854
rect 415102 204618 434546 204854
rect 434782 204618 434866 204854
rect 435102 204618 454546 204854
rect 454782 204618 454866 204854
rect 455102 204618 474546 204854
rect 474782 204618 474866 204854
rect 475102 204618 494546 204854
rect 494782 204618 494866 204854
rect 495102 204618 514546 204854
rect 514782 204618 514866 204854
rect 515102 204618 534546 204854
rect 534782 204618 534866 204854
rect 535102 204618 554546 204854
rect 554782 204618 554866 204854
rect 555102 204618 574546 204854
rect 574782 204618 574866 204854
rect 575102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 10826 201454
rect 11062 201218 11146 201454
rect 11382 201218 30826 201454
rect 31062 201218 31146 201454
rect 31382 201218 50826 201454
rect 51062 201218 51146 201454
rect 51382 201218 70826 201454
rect 71062 201218 71146 201454
rect 71382 201218 90826 201454
rect 91062 201218 91146 201454
rect 91382 201218 110826 201454
rect 111062 201218 111146 201454
rect 111382 201218 130826 201454
rect 131062 201218 131146 201454
rect 131382 201218 150826 201454
rect 151062 201218 151146 201454
rect 151382 201218 170826 201454
rect 171062 201218 171146 201454
rect 171382 201218 190826 201454
rect 191062 201218 191146 201454
rect 191382 201218 210826 201454
rect 211062 201218 211146 201454
rect 211382 201218 230826 201454
rect 231062 201218 231146 201454
rect 231382 201218 250826 201454
rect 251062 201218 251146 201454
rect 251382 201218 270826 201454
rect 271062 201218 271146 201454
rect 271382 201218 290826 201454
rect 291062 201218 291146 201454
rect 291382 201218 310826 201454
rect 311062 201218 311146 201454
rect 311382 201218 330826 201454
rect 331062 201218 331146 201454
rect 331382 201218 350826 201454
rect 351062 201218 351146 201454
rect 351382 201218 370826 201454
rect 371062 201218 371146 201454
rect 371382 201218 390826 201454
rect 391062 201218 391146 201454
rect 391382 201218 410826 201454
rect 411062 201218 411146 201454
rect 411382 201218 430826 201454
rect 431062 201218 431146 201454
rect 431382 201218 450826 201454
rect 451062 201218 451146 201454
rect 451382 201218 470826 201454
rect 471062 201218 471146 201454
rect 471382 201218 490826 201454
rect 491062 201218 491146 201454
rect 491382 201218 510826 201454
rect 511062 201218 511146 201454
rect 511382 201218 530826 201454
rect 531062 201218 531146 201454
rect 531382 201218 550826 201454
rect 551062 201218 551146 201454
rect 551382 201218 570826 201454
rect 571062 201218 571146 201454
rect 571382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 10826 201134
rect 11062 200898 11146 201134
rect 11382 200898 30826 201134
rect 31062 200898 31146 201134
rect 31382 200898 50826 201134
rect 51062 200898 51146 201134
rect 51382 200898 70826 201134
rect 71062 200898 71146 201134
rect 71382 200898 90826 201134
rect 91062 200898 91146 201134
rect 91382 200898 110826 201134
rect 111062 200898 111146 201134
rect 111382 200898 130826 201134
rect 131062 200898 131146 201134
rect 131382 200898 150826 201134
rect 151062 200898 151146 201134
rect 151382 200898 170826 201134
rect 171062 200898 171146 201134
rect 171382 200898 190826 201134
rect 191062 200898 191146 201134
rect 191382 200898 210826 201134
rect 211062 200898 211146 201134
rect 211382 200898 230826 201134
rect 231062 200898 231146 201134
rect 231382 200898 250826 201134
rect 251062 200898 251146 201134
rect 251382 200898 270826 201134
rect 271062 200898 271146 201134
rect 271382 200898 290826 201134
rect 291062 200898 291146 201134
rect 291382 200898 310826 201134
rect 311062 200898 311146 201134
rect 311382 200898 330826 201134
rect 331062 200898 331146 201134
rect 331382 200898 350826 201134
rect 351062 200898 351146 201134
rect 351382 200898 370826 201134
rect 371062 200898 371146 201134
rect 371382 200898 390826 201134
rect 391062 200898 391146 201134
rect 391382 200898 410826 201134
rect 411062 200898 411146 201134
rect 411382 200898 430826 201134
rect 431062 200898 431146 201134
rect 431382 200898 450826 201134
rect 451062 200898 451146 201134
rect 451382 200898 470826 201134
rect 471062 200898 471146 201134
rect 471382 200898 490826 201134
rect 491062 200898 491146 201134
rect 491382 200898 510826 201134
rect 511062 200898 511146 201134
rect 511382 200898 530826 201134
rect 531062 200898 531146 201134
rect 531382 200898 550826 201134
rect 551062 200898 551146 201134
rect 551382 200898 570826 201134
rect 571062 200898 571146 201134
rect 571382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 11986 194614
rect 12222 194378 12306 194614
rect 12542 194378 31986 194614
rect 32222 194378 32306 194614
rect 32542 194378 51986 194614
rect 52222 194378 52306 194614
rect 52542 194378 71986 194614
rect 72222 194378 72306 194614
rect 72542 194378 91986 194614
rect 92222 194378 92306 194614
rect 92542 194378 111986 194614
rect 112222 194378 112306 194614
rect 112542 194378 131986 194614
rect 132222 194378 132306 194614
rect 132542 194378 151986 194614
rect 152222 194378 152306 194614
rect 152542 194378 171986 194614
rect 172222 194378 172306 194614
rect 172542 194378 191986 194614
rect 192222 194378 192306 194614
rect 192542 194378 211986 194614
rect 212222 194378 212306 194614
rect 212542 194378 231986 194614
rect 232222 194378 232306 194614
rect 232542 194378 251986 194614
rect 252222 194378 252306 194614
rect 252542 194378 271986 194614
rect 272222 194378 272306 194614
rect 272542 194378 291986 194614
rect 292222 194378 292306 194614
rect 292542 194378 311986 194614
rect 312222 194378 312306 194614
rect 312542 194378 331986 194614
rect 332222 194378 332306 194614
rect 332542 194378 351986 194614
rect 352222 194378 352306 194614
rect 352542 194378 371986 194614
rect 372222 194378 372306 194614
rect 372542 194378 391986 194614
rect 392222 194378 392306 194614
rect 392542 194378 411986 194614
rect 412222 194378 412306 194614
rect 412542 194378 431986 194614
rect 432222 194378 432306 194614
rect 432542 194378 451986 194614
rect 452222 194378 452306 194614
rect 452542 194378 471986 194614
rect 472222 194378 472306 194614
rect 472542 194378 491986 194614
rect 492222 194378 492306 194614
rect 492542 194378 511986 194614
rect 512222 194378 512306 194614
rect 512542 194378 531986 194614
rect 532222 194378 532306 194614
rect 532542 194378 551986 194614
rect 552222 194378 552306 194614
rect 552542 194378 571986 194614
rect 572222 194378 572306 194614
rect 572542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 11986 194294
rect 12222 194058 12306 194294
rect 12542 194058 31986 194294
rect 32222 194058 32306 194294
rect 32542 194058 51986 194294
rect 52222 194058 52306 194294
rect 52542 194058 71986 194294
rect 72222 194058 72306 194294
rect 72542 194058 91986 194294
rect 92222 194058 92306 194294
rect 92542 194058 111986 194294
rect 112222 194058 112306 194294
rect 112542 194058 131986 194294
rect 132222 194058 132306 194294
rect 132542 194058 151986 194294
rect 152222 194058 152306 194294
rect 152542 194058 171986 194294
rect 172222 194058 172306 194294
rect 172542 194058 191986 194294
rect 192222 194058 192306 194294
rect 192542 194058 211986 194294
rect 212222 194058 212306 194294
rect 212542 194058 231986 194294
rect 232222 194058 232306 194294
rect 232542 194058 251986 194294
rect 252222 194058 252306 194294
rect 252542 194058 271986 194294
rect 272222 194058 272306 194294
rect 272542 194058 291986 194294
rect 292222 194058 292306 194294
rect 292542 194058 311986 194294
rect 312222 194058 312306 194294
rect 312542 194058 331986 194294
rect 332222 194058 332306 194294
rect 332542 194058 351986 194294
rect 352222 194058 352306 194294
rect 352542 194058 371986 194294
rect 372222 194058 372306 194294
rect 372542 194058 391986 194294
rect 392222 194058 392306 194294
rect 392542 194058 411986 194294
rect 412222 194058 412306 194294
rect 412542 194058 431986 194294
rect 432222 194058 432306 194294
rect 432542 194058 451986 194294
rect 452222 194058 452306 194294
rect 452542 194058 471986 194294
rect 472222 194058 472306 194294
rect 472542 194058 491986 194294
rect 492222 194058 492306 194294
rect 492542 194058 511986 194294
rect 512222 194058 512306 194294
rect 512542 194058 531986 194294
rect 532222 194058 532306 194294
rect 532542 194058 551986 194294
rect 552222 194058 552306 194294
rect 552542 194058 571986 194294
rect 572222 194058 572306 194294
rect 572542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 8266 190894
rect 8502 190658 8586 190894
rect 8822 190658 28266 190894
rect 28502 190658 28586 190894
rect 28822 190658 48266 190894
rect 48502 190658 48586 190894
rect 48822 190658 68266 190894
rect 68502 190658 68586 190894
rect 68822 190658 88266 190894
rect 88502 190658 88586 190894
rect 88822 190658 108266 190894
rect 108502 190658 108586 190894
rect 108822 190658 128266 190894
rect 128502 190658 128586 190894
rect 128822 190658 148266 190894
rect 148502 190658 148586 190894
rect 148822 190658 168266 190894
rect 168502 190658 168586 190894
rect 168822 190658 188266 190894
rect 188502 190658 188586 190894
rect 188822 190658 208266 190894
rect 208502 190658 208586 190894
rect 208822 190658 228266 190894
rect 228502 190658 228586 190894
rect 228822 190658 248266 190894
rect 248502 190658 248586 190894
rect 248822 190658 268266 190894
rect 268502 190658 268586 190894
rect 268822 190658 288266 190894
rect 288502 190658 288586 190894
rect 288822 190658 308266 190894
rect 308502 190658 308586 190894
rect 308822 190658 328266 190894
rect 328502 190658 328586 190894
rect 328822 190658 348266 190894
rect 348502 190658 348586 190894
rect 348822 190658 368266 190894
rect 368502 190658 368586 190894
rect 368822 190658 388266 190894
rect 388502 190658 388586 190894
rect 388822 190658 408266 190894
rect 408502 190658 408586 190894
rect 408822 190658 428266 190894
rect 428502 190658 428586 190894
rect 428822 190658 448266 190894
rect 448502 190658 448586 190894
rect 448822 190658 468266 190894
rect 468502 190658 468586 190894
rect 468822 190658 488266 190894
rect 488502 190658 488586 190894
rect 488822 190658 508266 190894
rect 508502 190658 508586 190894
rect 508822 190658 528266 190894
rect 528502 190658 528586 190894
rect 528822 190658 548266 190894
rect 548502 190658 548586 190894
rect 548822 190658 568266 190894
rect 568502 190658 568586 190894
rect 568822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 8266 190574
rect 8502 190338 8586 190574
rect 8822 190338 28266 190574
rect 28502 190338 28586 190574
rect 28822 190338 48266 190574
rect 48502 190338 48586 190574
rect 48822 190338 68266 190574
rect 68502 190338 68586 190574
rect 68822 190338 88266 190574
rect 88502 190338 88586 190574
rect 88822 190338 108266 190574
rect 108502 190338 108586 190574
rect 108822 190338 128266 190574
rect 128502 190338 128586 190574
rect 128822 190338 148266 190574
rect 148502 190338 148586 190574
rect 148822 190338 168266 190574
rect 168502 190338 168586 190574
rect 168822 190338 188266 190574
rect 188502 190338 188586 190574
rect 188822 190338 208266 190574
rect 208502 190338 208586 190574
rect 208822 190338 228266 190574
rect 228502 190338 228586 190574
rect 228822 190338 248266 190574
rect 248502 190338 248586 190574
rect 248822 190338 268266 190574
rect 268502 190338 268586 190574
rect 268822 190338 288266 190574
rect 288502 190338 288586 190574
rect 288822 190338 308266 190574
rect 308502 190338 308586 190574
rect 308822 190338 328266 190574
rect 328502 190338 328586 190574
rect 328822 190338 348266 190574
rect 348502 190338 348586 190574
rect 348822 190338 368266 190574
rect 368502 190338 368586 190574
rect 368822 190338 388266 190574
rect 388502 190338 388586 190574
rect 388822 190338 408266 190574
rect 408502 190338 408586 190574
rect 408822 190338 428266 190574
rect 428502 190338 428586 190574
rect 428822 190338 448266 190574
rect 448502 190338 448586 190574
rect 448822 190338 468266 190574
rect 468502 190338 468586 190574
rect 468822 190338 488266 190574
rect 488502 190338 488586 190574
rect 488822 190338 508266 190574
rect 508502 190338 508586 190574
rect 508822 190338 528266 190574
rect 528502 190338 528586 190574
rect 528822 190338 548266 190574
rect 548502 190338 548586 190574
rect 548822 190338 568266 190574
rect 568502 190338 568586 190574
rect 568822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 4546 187174
rect 4782 186938 4866 187174
rect 5102 186938 24546 187174
rect 24782 186938 24866 187174
rect 25102 186938 44546 187174
rect 44782 186938 44866 187174
rect 45102 186938 64546 187174
rect 64782 186938 64866 187174
rect 65102 186938 84546 187174
rect 84782 186938 84866 187174
rect 85102 186938 104546 187174
rect 104782 186938 104866 187174
rect 105102 186938 124546 187174
rect 124782 186938 124866 187174
rect 125102 186938 144546 187174
rect 144782 186938 144866 187174
rect 145102 186938 164546 187174
rect 164782 186938 164866 187174
rect 165102 186938 184546 187174
rect 184782 186938 184866 187174
rect 185102 186938 204546 187174
rect 204782 186938 204866 187174
rect 205102 186938 224546 187174
rect 224782 186938 224866 187174
rect 225102 186938 244546 187174
rect 244782 186938 244866 187174
rect 245102 186938 264546 187174
rect 264782 186938 264866 187174
rect 265102 186938 284546 187174
rect 284782 186938 284866 187174
rect 285102 186938 304546 187174
rect 304782 186938 304866 187174
rect 305102 186938 324546 187174
rect 324782 186938 324866 187174
rect 325102 186938 344546 187174
rect 344782 186938 344866 187174
rect 345102 186938 364546 187174
rect 364782 186938 364866 187174
rect 365102 186938 384546 187174
rect 384782 186938 384866 187174
rect 385102 186938 404546 187174
rect 404782 186938 404866 187174
rect 405102 186938 424546 187174
rect 424782 186938 424866 187174
rect 425102 186938 444546 187174
rect 444782 186938 444866 187174
rect 445102 186938 464546 187174
rect 464782 186938 464866 187174
rect 465102 186938 484546 187174
rect 484782 186938 484866 187174
rect 485102 186938 504546 187174
rect 504782 186938 504866 187174
rect 505102 186938 524546 187174
rect 524782 186938 524866 187174
rect 525102 186938 544546 187174
rect 544782 186938 544866 187174
rect 545102 186938 564546 187174
rect 564782 186938 564866 187174
rect 565102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 4546 186854
rect 4782 186618 4866 186854
rect 5102 186618 24546 186854
rect 24782 186618 24866 186854
rect 25102 186618 44546 186854
rect 44782 186618 44866 186854
rect 45102 186618 64546 186854
rect 64782 186618 64866 186854
rect 65102 186618 84546 186854
rect 84782 186618 84866 186854
rect 85102 186618 104546 186854
rect 104782 186618 104866 186854
rect 105102 186618 124546 186854
rect 124782 186618 124866 186854
rect 125102 186618 144546 186854
rect 144782 186618 144866 186854
rect 145102 186618 164546 186854
rect 164782 186618 164866 186854
rect 165102 186618 184546 186854
rect 184782 186618 184866 186854
rect 185102 186618 204546 186854
rect 204782 186618 204866 186854
rect 205102 186618 224546 186854
rect 224782 186618 224866 186854
rect 225102 186618 244546 186854
rect 244782 186618 244866 186854
rect 245102 186618 264546 186854
rect 264782 186618 264866 186854
rect 265102 186618 284546 186854
rect 284782 186618 284866 186854
rect 285102 186618 304546 186854
rect 304782 186618 304866 186854
rect 305102 186618 324546 186854
rect 324782 186618 324866 186854
rect 325102 186618 344546 186854
rect 344782 186618 344866 186854
rect 345102 186618 364546 186854
rect 364782 186618 364866 186854
rect 365102 186618 384546 186854
rect 384782 186618 384866 186854
rect 385102 186618 404546 186854
rect 404782 186618 404866 186854
rect 405102 186618 424546 186854
rect 424782 186618 424866 186854
rect 425102 186618 444546 186854
rect 444782 186618 444866 186854
rect 445102 186618 464546 186854
rect 464782 186618 464866 186854
rect 465102 186618 484546 186854
rect 484782 186618 484866 186854
rect 485102 186618 504546 186854
rect 504782 186618 504866 186854
rect 505102 186618 524546 186854
rect 524782 186618 524866 186854
rect 525102 186618 544546 186854
rect 544782 186618 544866 186854
rect 545102 186618 564546 186854
rect 564782 186618 564866 186854
rect 565102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 826 183454
rect 1062 183218 1146 183454
rect 1382 183218 20826 183454
rect 21062 183218 21146 183454
rect 21382 183218 40826 183454
rect 41062 183218 41146 183454
rect 41382 183218 60826 183454
rect 61062 183218 61146 183454
rect 61382 183218 80826 183454
rect 81062 183218 81146 183454
rect 81382 183218 100826 183454
rect 101062 183218 101146 183454
rect 101382 183218 120826 183454
rect 121062 183218 121146 183454
rect 121382 183218 140826 183454
rect 141062 183218 141146 183454
rect 141382 183218 160826 183454
rect 161062 183218 161146 183454
rect 161382 183218 180826 183454
rect 181062 183218 181146 183454
rect 181382 183218 200826 183454
rect 201062 183218 201146 183454
rect 201382 183218 220826 183454
rect 221062 183218 221146 183454
rect 221382 183218 240826 183454
rect 241062 183218 241146 183454
rect 241382 183218 260826 183454
rect 261062 183218 261146 183454
rect 261382 183218 280826 183454
rect 281062 183218 281146 183454
rect 281382 183218 300826 183454
rect 301062 183218 301146 183454
rect 301382 183218 320826 183454
rect 321062 183218 321146 183454
rect 321382 183218 340826 183454
rect 341062 183218 341146 183454
rect 341382 183218 360826 183454
rect 361062 183218 361146 183454
rect 361382 183218 380826 183454
rect 381062 183218 381146 183454
rect 381382 183218 400826 183454
rect 401062 183218 401146 183454
rect 401382 183218 420826 183454
rect 421062 183218 421146 183454
rect 421382 183218 440826 183454
rect 441062 183218 441146 183454
rect 441382 183218 460826 183454
rect 461062 183218 461146 183454
rect 461382 183218 480826 183454
rect 481062 183218 481146 183454
rect 481382 183218 500826 183454
rect 501062 183218 501146 183454
rect 501382 183218 520826 183454
rect 521062 183218 521146 183454
rect 521382 183218 540826 183454
rect 541062 183218 541146 183454
rect 541382 183218 560826 183454
rect 561062 183218 561146 183454
rect 561382 183218 580826 183454
rect 581062 183218 581146 183454
rect 581382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 826 183134
rect 1062 182898 1146 183134
rect 1382 182898 20826 183134
rect 21062 182898 21146 183134
rect 21382 182898 40826 183134
rect 41062 182898 41146 183134
rect 41382 182898 60826 183134
rect 61062 182898 61146 183134
rect 61382 182898 80826 183134
rect 81062 182898 81146 183134
rect 81382 182898 100826 183134
rect 101062 182898 101146 183134
rect 101382 182898 120826 183134
rect 121062 182898 121146 183134
rect 121382 182898 140826 183134
rect 141062 182898 141146 183134
rect 141382 182898 160826 183134
rect 161062 182898 161146 183134
rect 161382 182898 180826 183134
rect 181062 182898 181146 183134
rect 181382 182898 200826 183134
rect 201062 182898 201146 183134
rect 201382 182898 220826 183134
rect 221062 182898 221146 183134
rect 221382 182898 240826 183134
rect 241062 182898 241146 183134
rect 241382 182898 260826 183134
rect 261062 182898 261146 183134
rect 261382 182898 280826 183134
rect 281062 182898 281146 183134
rect 281382 182898 300826 183134
rect 301062 182898 301146 183134
rect 301382 182898 320826 183134
rect 321062 182898 321146 183134
rect 321382 182898 340826 183134
rect 341062 182898 341146 183134
rect 341382 182898 360826 183134
rect 361062 182898 361146 183134
rect 361382 182898 380826 183134
rect 381062 182898 381146 183134
rect 381382 182898 400826 183134
rect 401062 182898 401146 183134
rect 401382 182898 420826 183134
rect 421062 182898 421146 183134
rect 421382 182898 440826 183134
rect 441062 182898 441146 183134
rect 441382 182898 460826 183134
rect 461062 182898 461146 183134
rect 461382 182898 480826 183134
rect 481062 182898 481146 183134
rect 481382 182898 500826 183134
rect 501062 182898 501146 183134
rect 501382 182898 520826 183134
rect 521062 182898 521146 183134
rect 521382 182898 540826 183134
rect 541062 182898 541146 183134
rect 541382 182898 560826 183134
rect 561062 182898 561146 183134
rect 561382 182898 580826 183134
rect 581062 182898 581146 183134
rect 581382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 21986 176614
rect 22222 176378 22306 176614
rect 22542 176378 41986 176614
rect 42222 176378 42306 176614
rect 42542 176378 61986 176614
rect 62222 176378 62306 176614
rect 62542 176378 81986 176614
rect 82222 176378 82306 176614
rect 82542 176378 101986 176614
rect 102222 176378 102306 176614
rect 102542 176378 121986 176614
rect 122222 176378 122306 176614
rect 122542 176378 141986 176614
rect 142222 176378 142306 176614
rect 142542 176378 161986 176614
rect 162222 176378 162306 176614
rect 162542 176378 181986 176614
rect 182222 176378 182306 176614
rect 182542 176378 201986 176614
rect 202222 176378 202306 176614
rect 202542 176378 221986 176614
rect 222222 176378 222306 176614
rect 222542 176378 241986 176614
rect 242222 176378 242306 176614
rect 242542 176378 261986 176614
rect 262222 176378 262306 176614
rect 262542 176378 281986 176614
rect 282222 176378 282306 176614
rect 282542 176378 301986 176614
rect 302222 176378 302306 176614
rect 302542 176378 321986 176614
rect 322222 176378 322306 176614
rect 322542 176378 341986 176614
rect 342222 176378 342306 176614
rect 342542 176378 361986 176614
rect 362222 176378 362306 176614
rect 362542 176378 381986 176614
rect 382222 176378 382306 176614
rect 382542 176378 401986 176614
rect 402222 176378 402306 176614
rect 402542 176378 421986 176614
rect 422222 176378 422306 176614
rect 422542 176378 441986 176614
rect 442222 176378 442306 176614
rect 442542 176378 461986 176614
rect 462222 176378 462306 176614
rect 462542 176378 481986 176614
rect 482222 176378 482306 176614
rect 482542 176378 501986 176614
rect 502222 176378 502306 176614
rect 502542 176378 521986 176614
rect 522222 176378 522306 176614
rect 522542 176378 541986 176614
rect 542222 176378 542306 176614
rect 542542 176378 561986 176614
rect 562222 176378 562306 176614
rect 562542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 21986 176294
rect 22222 176058 22306 176294
rect 22542 176058 41986 176294
rect 42222 176058 42306 176294
rect 42542 176058 61986 176294
rect 62222 176058 62306 176294
rect 62542 176058 81986 176294
rect 82222 176058 82306 176294
rect 82542 176058 101986 176294
rect 102222 176058 102306 176294
rect 102542 176058 121986 176294
rect 122222 176058 122306 176294
rect 122542 176058 141986 176294
rect 142222 176058 142306 176294
rect 142542 176058 161986 176294
rect 162222 176058 162306 176294
rect 162542 176058 181986 176294
rect 182222 176058 182306 176294
rect 182542 176058 201986 176294
rect 202222 176058 202306 176294
rect 202542 176058 221986 176294
rect 222222 176058 222306 176294
rect 222542 176058 241986 176294
rect 242222 176058 242306 176294
rect 242542 176058 261986 176294
rect 262222 176058 262306 176294
rect 262542 176058 281986 176294
rect 282222 176058 282306 176294
rect 282542 176058 301986 176294
rect 302222 176058 302306 176294
rect 302542 176058 321986 176294
rect 322222 176058 322306 176294
rect 322542 176058 341986 176294
rect 342222 176058 342306 176294
rect 342542 176058 361986 176294
rect 362222 176058 362306 176294
rect 362542 176058 381986 176294
rect 382222 176058 382306 176294
rect 382542 176058 401986 176294
rect 402222 176058 402306 176294
rect 402542 176058 421986 176294
rect 422222 176058 422306 176294
rect 422542 176058 441986 176294
rect 442222 176058 442306 176294
rect 442542 176058 461986 176294
rect 462222 176058 462306 176294
rect 462542 176058 481986 176294
rect 482222 176058 482306 176294
rect 482542 176058 501986 176294
rect 502222 176058 502306 176294
rect 502542 176058 521986 176294
rect 522222 176058 522306 176294
rect 522542 176058 541986 176294
rect 542222 176058 542306 176294
rect 542542 176058 561986 176294
rect 562222 176058 562306 176294
rect 562542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 18266 172894
rect 18502 172658 18586 172894
rect 18822 172658 38266 172894
rect 38502 172658 38586 172894
rect 38822 172658 58266 172894
rect 58502 172658 58586 172894
rect 58822 172658 78266 172894
rect 78502 172658 78586 172894
rect 78822 172658 98266 172894
rect 98502 172658 98586 172894
rect 98822 172658 118266 172894
rect 118502 172658 118586 172894
rect 118822 172658 138266 172894
rect 138502 172658 138586 172894
rect 138822 172658 158266 172894
rect 158502 172658 158586 172894
rect 158822 172658 178266 172894
rect 178502 172658 178586 172894
rect 178822 172658 198266 172894
rect 198502 172658 198586 172894
rect 198822 172658 218266 172894
rect 218502 172658 218586 172894
rect 218822 172658 238266 172894
rect 238502 172658 238586 172894
rect 238822 172658 258266 172894
rect 258502 172658 258586 172894
rect 258822 172658 278266 172894
rect 278502 172658 278586 172894
rect 278822 172658 298266 172894
rect 298502 172658 298586 172894
rect 298822 172658 318266 172894
rect 318502 172658 318586 172894
rect 318822 172658 338266 172894
rect 338502 172658 338586 172894
rect 338822 172658 358266 172894
rect 358502 172658 358586 172894
rect 358822 172658 378266 172894
rect 378502 172658 378586 172894
rect 378822 172658 398266 172894
rect 398502 172658 398586 172894
rect 398822 172658 418266 172894
rect 418502 172658 418586 172894
rect 418822 172658 438266 172894
rect 438502 172658 438586 172894
rect 438822 172658 458266 172894
rect 458502 172658 458586 172894
rect 458822 172658 478266 172894
rect 478502 172658 478586 172894
rect 478822 172658 498266 172894
rect 498502 172658 498586 172894
rect 498822 172658 518266 172894
rect 518502 172658 518586 172894
rect 518822 172658 538266 172894
rect 538502 172658 538586 172894
rect 538822 172658 558266 172894
rect 558502 172658 558586 172894
rect 558822 172658 578266 172894
rect 578502 172658 578586 172894
rect 578822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 18266 172574
rect 18502 172338 18586 172574
rect 18822 172338 38266 172574
rect 38502 172338 38586 172574
rect 38822 172338 58266 172574
rect 58502 172338 58586 172574
rect 58822 172338 78266 172574
rect 78502 172338 78586 172574
rect 78822 172338 98266 172574
rect 98502 172338 98586 172574
rect 98822 172338 118266 172574
rect 118502 172338 118586 172574
rect 118822 172338 138266 172574
rect 138502 172338 138586 172574
rect 138822 172338 158266 172574
rect 158502 172338 158586 172574
rect 158822 172338 178266 172574
rect 178502 172338 178586 172574
rect 178822 172338 198266 172574
rect 198502 172338 198586 172574
rect 198822 172338 218266 172574
rect 218502 172338 218586 172574
rect 218822 172338 238266 172574
rect 238502 172338 238586 172574
rect 238822 172338 258266 172574
rect 258502 172338 258586 172574
rect 258822 172338 278266 172574
rect 278502 172338 278586 172574
rect 278822 172338 298266 172574
rect 298502 172338 298586 172574
rect 298822 172338 318266 172574
rect 318502 172338 318586 172574
rect 318822 172338 338266 172574
rect 338502 172338 338586 172574
rect 338822 172338 358266 172574
rect 358502 172338 358586 172574
rect 358822 172338 378266 172574
rect 378502 172338 378586 172574
rect 378822 172338 398266 172574
rect 398502 172338 398586 172574
rect 398822 172338 418266 172574
rect 418502 172338 418586 172574
rect 418822 172338 438266 172574
rect 438502 172338 438586 172574
rect 438822 172338 458266 172574
rect 458502 172338 458586 172574
rect 458822 172338 478266 172574
rect 478502 172338 478586 172574
rect 478822 172338 498266 172574
rect 498502 172338 498586 172574
rect 498822 172338 518266 172574
rect 518502 172338 518586 172574
rect 518822 172338 538266 172574
rect 538502 172338 538586 172574
rect 538822 172338 558266 172574
rect 558502 172338 558586 172574
rect 558822 172338 578266 172574
rect 578502 172338 578586 172574
rect 578822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 14546 169174
rect 14782 168938 14866 169174
rect 15102 168938 34546 169174
rect 34782 168938 34866 169174
rect 35102 168938 54546 169174
rect 54782 168938 54866 169174
rect 55102 168938 74546 169174
rect 74782 168938 74866 169174
rect 75102 168938 94546 169174
rect 94782 168938 94866 169174
rect 95102 168938 114546 169174
rect 114782 168938 114866 169174
rect 115102 168938 134546 169174
rect 134782 168938 134866 169174
rect 135102 168938 154546 169174
rect 154782 168938 154866 169174
rect 155102 168938 174546 169174
rect 174782 168938 174866 169174
rect 175102 168938 194546 169174
rect 194782 168938 194866 169174
rect 195102 168938 214546 169174
rect 214782 168938 214866 169174
rect 215102 168938 234546 169174
rect 234782 168938 234866 169174
rect 235102 168938 254546 169174
rect 254782 168938 254866 169174
rect 255102 168938 274546 169174
rect 274782 168938 274866 169174
rect 275102 168938 294546 169174
rect 294782 168938 294866 169174
rect 295102 168938 314546 169174
rect 314782 168938 314866 169174
rect 315102 168938 334546 169174
rect 334782 168938 334866 169174
rect 335102 168938 354546 169174
rect 354782 168938 354866 169174
rect 355102 168938 374546 169174
rect 374782 168938 374866 169174
rect 375102 168938 394546 169174
rect 394782 168938 394866 169174
rect 395102 168938 414546 169174
rect 414782 168938 414866 169174
rect 415102 168938 434546 169174
rect 434782 168938 434866 169174
rect 435102 168938 454546 169174
rect 454782 168938 454866 169174
rect 455102 168938 474546 169174
rect 474782 168938 474866 169174
rect 475102 168938 494546 169174
rect 494782 168938 494866 169174
rect 495102 168938 514546 169174
rect 514782 168938 514866 169174
rect 515102 168938 534546 169174
rect 534782 168938 534866 169174
rect 535102 168938 554546 169174
rect 554782 168938 554866 169174
rect 555102 168938 574546 169174
rect 574782 168938 574866 169174
rect 575102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 14546 168854
rect 14782 168618 14866 168854
rect 15102 168618 34546 168854
rect 34782 168618 34866 168854
rect 35102 168618 54546 168854
rect 54782 168618 54866 168854
rect 55102 168618 74546 168854
rect 74782 168618 74866 168854
rect 75102 168618 94546 168854
rect 94782 168618 94866 168854
rect 95102 168618 114546 168854
rect 114782 168618 114866 168854
rect 115102 168618 134546 168854
rect 134782 168618 134866 168854
rect 135102 168618 154546 168854
rect 154782 168618 154866 168854
rect 155102 168618 174546 168854
rect 174782 168618 174866 168854
rect 175102 168618 194546 168854
rect 194782 168618 194866 168854
rect 195102 168618 214546 168854
rect 214782 168618 214866 168854
rect 215102 168618 234546 168854
rect 234782 168618 234866 168854
rect 235102 168618 254546 168854
rect 254782 168618 254866 168854
rect 255102 168618 274546 168854
rect 274782 168618 274866 168854
rect 275102 168618 294546 168854
rect 294782 168618 294866 168854
rect 295102 168618 314546 168854
rect 314782 168618 314866 168854
rect 315102 168618 334546 168854
rect 334782 168618 334866 168854
rect 335102 168618 354546 168854
rect 354782 168618 354866 168854
rect 355102 168618 374546 168854
rect 374782 168618 374866 168854
rect 375102 168618 394546 168854
rect 394782 168618 394866 168854
rect 395102 168618 414546 168854
rect 414782 168618 414866 168854
rect 415102 168618 434546 168854
rect 434782 168618 434866 168854
rect 435102 168618 454546 168854
rect 454782 168618 454866 168854
rect 455102 168618 474546 168854
rect 474782 168618 474866 168854
rect 475102 168618 494546 168854
rect 494782 168618 494866 168854
rect 495102 168618 514546 168854
rect 514782 168618 514866 168854
rect 515102 168618 534546 168854
rect 534782 168618 534866 168854
rect 535102 168618 554546 168854
rect 554782 168618 554866 168854
rect 555102 168618 574546 168854
rect 574782 168618 574866 168854
rect 575102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 10826 165454
rect 11062 165218 11146 165454
rect 11382 165218 30826 165454
rect 31062 165218 31146 165454
rect 31382 165218 50826 165454
rect 51062 165218 51146 165454
rect 51382 165218 70826 165454
rect 71062 165218 71146 165454
rect 71382 165218 90826 165454
rect 91062 165218 91146 165454
rect 91382 165218 110826 165454
rect 111062 165218 111146 165454
rect 111382 165218 130826 165454
rect 131062 165218 131146 165454
rect 131382 165218 150826 165454
rect 151062 165218 151146 165454
rect 151382 165218 170826 165454
rect 171062 165218 171146 165454
rect 171382 165218 190826 165454
rect 191062 165218 191146 165454
rect 191382 165218 210826 165454
rect 211062 165218 211146 165454
rect 211382 165218 230826 165454
rect 231062 165218 231146 165454
rect 231382 165218 250826 165454
rect 251062 165218 251146 165454
rect 251382 165218 270826 165454
rect 271062 165218 271146 165454
rect 271382 165218 290826 165454
rect 291062 165218 291146 165454
rect 291382 165218 310826 165454
rect 311062 165218 311146 165454
rect 311382 165218 330826 165454
rect 331062 165218 331146 165454
rect 331382 165218 350826 165454
rect 351062 165218 351146 165454
rect 351382 165218 370826 165454
rect 371062 165218 371146 165454
rect 371382 165218 390826 165454
rect 391062 165218 391146 165454
rect 391382 165218 410826 165454
rect 411062 165218 411146 165454
rect 411382 165218 430826 165454
rect 431062 165218 431146 165454
rect 431382 165218 450826 165454
rect 451062 165218 451146 165454
rect 451382 165218 470826 165454
rect 471062 165218 471146 165454
rect 471382 165218 490826 165454
rect 491062 165218 491146 165454
rect 491382 165218 510826 165454
rect 511062 165218 511146 165454
rect 511382 165218 530826 165454
rect 531062 165218 531146 165454
rect 531382 165218 550826 165454
rect 551062 165218 551146 165454
rect 551382 165218 570826 165454
rect 571062 165218 571146 165454
rect 571382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 10826 165134
rect 11062 164898 11146 165134
rect 11382 164898 30826 165134
rect 31062 164898 31146 165134
rect 31382 164898 50826 165134
rect 51062 164898 51146 165134
rect 51382 164898 70826 165134
rect 71062 164898 71146 165134
rect 71382 164898 90826 165134
rect 91062 164898 91146 165134
rect 91382 164898 110826 165134
rect 111062 164898 111146 165134
rect 111382 164898 130826 165134
rect 131062 164898 131146 165134
rect 131382 164898 150826 165134
rect 151062 164898 151146 165134
rect 151382 164898 170826 165134
rect 171062 164898 171146 165134
rect 171382 164898 190826 165134
rect 191062 164898 191146 165134
rect 191382 164898 210826 165134
rect 211062 164898 211146 165134
rect 211382 164898 230826 165134
rect 231062 164898 231146 165134
rect 231382 164898 250826 165134
rect 251062 164898 251146 165134
rect 251382 164898 270826 165134
rect 271062 164898 271146 165134
rect 271382 164898 290826 165134
rect 291062 164898 291146 165134
rect 291382 164898 310826 165134
rect 311062 164898 311146 165134
rect 311382 164898 330826 165134
rect 331062 164898 331146 165134
rect 331382 164898 350826 165134
rect 351062 164898 351146 165134
rect 351382 164898 370826 165134
rect 371062 164898 371146 165134
rect 371382 164898 390826 165134
rect 391062 164898 391146 165134
rect 391382 164898 410826 165134
rect 411062 164898 411146 165134
rect 411382 164898 430826 165134
rect 431062 164898 431146 165134
rect 431382 164898 450826 165134
rect 451062 164898 451146 165134
rect 451382 164898 470826 165134
rect 471062 164898 471146 165134
rect 471382 164898 490826 165134
rect 491062 164898 491146 165134
rect 491382 164898 510826 165134
rect 511062 164898 511146 165134
rect 511382 164898 530826 165134
rect 531062 164898 531146 165134
rect 531382 164898 550826 165134
rect 551062 164898 551146 165134
rect 551382 164898 570826 165134
rect 571062 164898 571146 165134
rect 571382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 11986 158614
rect 12222 158378 12306 158614
rect 12542 158378 31986 158614
rect 32222 158378 32306 158614
rect 32542 158378 51986 158614
rect 52222 158378 52306 158614
rect 52542 158378 71986 158614
rect 72222 158378 72306 158614
rect 72542 158378 91986 158614
rect 92222 158378 92306 158614
rect 92542 158378 111986 158614
rect 112222 158378 112306 158614
rect 112542 158378 131986 158614
rect 132222 158378 132306 158614
rect 132542 158378 151986 158614
rect 152222 158378 152306 158614
rect 152542 158378 171986 158614
rect 172222 158378 172306 158614
rect 172542 158378 191986 158614
rect 192222 158378 192306 158614
rect 192542 158378 211986 158614
rect 212222 158378 212306 158614
rect 212542 158378 231986 158614
rect 232222 158378 232306 158614
rect 232542 158378 251986 158614
rect 252222 158378 252306 158614
rect 252542 158378 271986 158614
rect 272222 158378 272306 158614
rect 272542 158378 291986 158614
rect 292222 158378 292306 158614
rect 292542 158378 311986 158614
rect 312222 158378 312306 158614
rect 312542 158378 331986 158614
rect 332222 158378 332306 158614
rect 332542 158378 351986 158614
rect 352222 158378 352306 158614
rect 352542 158378 371986 158614
rect 372222 158378 372306 158614
rect 372542 158378 391986 158614
rect 392222 158378 392306 158614
rect 392542 158378 411986 158614
rect 412222 158378 412306 158614
rect 412542 158378 431986 158614
rect 432222 158378 432306 158614
rect 432542 158378 451986 158614
rect 452222 158378 452306 158614
rect 452542 158378 471986 158614
rect 472222 158378 472306 158614
rect 472542 158378 491986 158614
rect 492222 158378 492306 158614
rect 492542 158378 511986 158614
rect 512222 158378 512306 158614
rect 512542 158378 531986 158614
rect 532222 158378 532306 158614
rect 532542 158378 551986 158614
rect 552222 158378 552306 158614
rect 552542 158378 571986 158614
rect 572222 158378 572306 158614
rect 572542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 11986 158294
rect 12222 158058 12306 158294
rect 12542 158058 31986 158294
rect 32222 158058 32306 158294
rect 32542 158058 51986 158294
rect 52222 158058 52306 158294
rect 52542 158058 71986 158294
rect 72222 158058 72306 158294
rect 72542 158058 91986 158294
rect 92222 158058 92306 158294
rect 92542 158058 111986 158294
rect 112222 158058 112306 158294
rect 112542 158058 131986 158294
rect 132222 158058 132306 158294
rect 132542 158058 151986 158294
rect 152222 158058 152306 158294
rect 152542 158058 171986 158294
rect 172222 158058 172306 158294
rect 172542 158058 191986 158294
rect 192222 158058 192306 158294
rect 192542 158058 211986 158294
rect 212222 158058 212306 158294
rect 212542 158058 231986 158294
rect 232222 158058 232306 158294
rect 232542 158058 251986 158294
rect 252222 158058 252306 158294
rect 252542 158058 271986 158294
rect 272222 158058 272306 158294
rect 272542 158058 291986 158294
rect 292222 158058 292306 158294
rect 292542 158058 311986 158294
rect 312222 158058 312306 158294
rect 312542 158058 331986 158294
rect 332222 158058 332306 158294
rect 332542 158058 351986 158294
rect 352222 158058 352306 158294
rect 352542 158058 371986 158294
rect 372222 158058 372306 158294
rect 372542 158058 391986 158294
rect 392222 158058 392306 158294
rect 392542 158058 411986 158294
rect 412222 158058 412306 158294
rect 412542 158058 431986 158294
rect 432222 158058 432306 158294
rect 432542 158058 451986 158294
rect 452222 158058 452306 158294
rect 452542 158058 471986 158294
rect 472222 158058 472306 158294
rect 472542 158058 491986 158294
rect 492222 158058 492306 158294
rect 492542 158058 511986 158294
rect 512222 158058 512306 158294
rect 512542 158058 531986 158294
rect 532222 158058 532306 158294
rect 532542 158058 551986 158294
rect 552222 158058 552306 158294
rect 552542 158058 571986 158294
rect 572222 158058 572306 158294
rect 572542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 8266 154894
rect 8502 154658 8586 154894
rect 8822 154658 28266 154894
rect 28502 154658 28586 154894
rect 28822 154658 48266 154894
rect 48502 154658 48586 154894
rect 48822 154658 68266 154894
rect 68502 154658 68586 154894
rect 68822 154658 88266 154894
rect 88502 154658 88586 154894
rect 88822 154658 108266 154894
rect 108502 154658 108586 154894
rect 108822 154658 128266 154894
rect 128502 154658 128586 154894
rect 128822 154658 148266 154894
rect 148502 154658 148586 154894
rect 148822 154658 168266 154894
rect 168502 154658 168586 154894
rect 168822 154658 188266 154894
rect 188502 154658 188586 154894
rect 188822 154658 208266 154894
rect 208502 154658 208586 154894
rect 208822 154658 228266 154894
rect 228502 154658 228586 154894
rect 228822 154658 248266 154894
rect 248502 154658 248586 154894
rect 248822 154658 268266 154894
rect 268502 154658 268586 154894
rect 268822 154658 288266 154894
rect 288502 154658 288586 154894
rect 288822 154658 308266 154894
rect 308502 154658 308586 154894
rect 308822 154658 328266 154894
rect 328502 154658 328586 154894
rect 328822 154658 348266 154894
rect 348502 154658 348586 154894
rect 348822 154658 368266 154894
rect 368502 154658 368586 154894
rect 368822 154658 388266 154894
rect 388502 154658 388586 154894
rect 388822 154658 408266 154894
rect 408502 154658 408586 154894
rect 408822 154658 428266 154894
rect 428502 154658 428586 154894
rect 428822 154658 448266 154894
rect 448502 154658 448586 154894
rect 448822 154658 468266 154894
rect 468502 154658 468586 154894
rect 468822 154658 488266 154894
rect 488502 154658 488586 154894
rect 488822 154658 508266 154894
rect 508502 154658 508586 154894
rect 508822 154658 528266 154894
rect 528502 154658 528586 154894
rect 528822 154658 548266 154894
rect 548502 154658 548586 154894
rect 548822 154658 568266 154894
rect 568502 154658 568586 154894
rect 568822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 8266 154574
rect 8502 154338 8586 154574
rect 8822 154338 28266 154574
rect 28502 154338 28586 154574
rect 28822 154338 48266 154574
rect 48502 154338 48586 154574
rect 48822 154338 68266 154574
rect 68502 154338 68586 154574
rect 68822 154338 88266 154574
rect 88502 154338 88586 154574
rect 88822 154338 108266 154574
rect 108502 154338 108586 154574
rect 108822 154338 128266 154574
rect 128502 154338 128586 154574
rect 128822 154338 148266 154574
rect 148502 154338 148586 154574
rect 148822 154338 168266 154574
rect 168502 154338 168586 154574
rect 168822 154338 188266 154574
rect 188502 154338 188586 154574
rect 188822 154338 208266 154574
rect 208502 154338 208586 154574
rect 208822 154338 228266 154574
rect 228502 154338 228586 154574
rect 228822 154338 248266 154574
rect 248502 154338 248586 154574
rect 248822 154338 268266 154574
rect 268502 154338 268586 154574
rect 268822 154338 288266 154574
rect 288502 154338 288586 154574
rect 288822 154338 308266 154574
rect 308502 154338 308586 154574
rect 308822 154338 328266 154574
rect 328502 154338 328586 154574
rect 328822 154338 348266 154574
rect 348502 154338 348586 154574
rect 348822 154338 368266 154574
rect 368502 154338 368586 154574
rect 368822 154338 388266 154574
rect 388502 154338 388586 154574
rect 388822 154338 408266 154574
rect 408502 154338 408586 154574
rect 408822 154338 428266 154574
rect 428502 154338 428586 154574
rect 428822 154338 448266 154574
rect 448502 154338 448586 154574
rect 448822 154338 468266 154574
rect 468502 154338 468586 154574
rect 468822 154338 488266 154574
rect 488502 154338 488586 154574
rect 488822 154338 508266 154574
rect 508502 154338 508586 154574
rect 508822 154338 528266 154574
rect 528502 154338 528586 154574
rect 528822 154338 548266 154574
rect 548502 154338 548586 154574
rect 548822 154338 568266 154574
rect 568502 154338 568586 154574
rect 568822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 4546 151174
rect 4782 150938 4866 151174
rect 5102 150938 24546 151174
rect 24782 150938 24866 151174
rect 25102 150938 44546 151174
rect 44782 150938 44866 151174
rect 45102 150938 64546 151174
rect 64782 150938 64866 151174
rect 65102 150938 84546 151174
rect 84782 150938 84866 151174
rect 85102 150938 104546 151174
rect 104782 150938 104866 151174
rect 105102 150938 124546 151174
rect 124782 150938 124866 151174
rect 125102 150938 144546 151174
rect 144782 150938 144866 151174
rect 145102 150938 164546 151174
rect 164782 150938 164866 151174
rect 165102 150938 184546 151174
rect 184782 150938 184866 151174
rect 185102 150938 204546 151174
rect 204782 150938 204866 151174
rect 205102 150938 224546 151174
rect 224782 150938 224866 151174
rect 225102 150938 244546 151174
rect 244782 150938 244866 151174
rect 245102 150938 264546 151174
rect 264782 150938 264866 151174
rect 265102 150938 284546 151174
rect 284782 150938 284866 151174
rect 285102 150938 304546 151174
rect 304782 150938 304866 151174
rect 305102 150938 324546 151174
rect 324782 150938 324866 151174
rect 325102 150938 344546 151174
rect 344782 150938 344866 151174
rect 345102 150938 364546 151174
rect 364782 150938 364866 151174
rect 365102 150938 384546 151174
rect 384782 150938 384866 151174
rect 385102 150938 404546 151174
rect 404782 150938 404866 151174
rect 405102 150938 424546 151174
rect 424782 150938 424866 151174
rect 425102 150938 444546 151174
rect 444782 150938 444866 151174
rect 445102 150938 464546 151174
rect 464782 150938 464866 151174
rect 465102 150938 484546 151174
rect 484782 150938 484866 151174
rect 485102 150938 504546 151174
rect 504782 150938 504866 151174
rect 505102 150938 524546 151174
rect 524782 150938 524866 151174
rect 525102 150938 544546 151174
rect 544782 150938 544866 151174
rect 545102 150938 564546 151174
rect 564782 150938 564866 151174
rect 565102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 4546 150854
rect 4782 150618 4866 150854
rect 5102 150618 24546 150854
rect 24782 150618 24866 150854
rect 25102 150618 44546 150854
rect 44782 150618 44866 150854
rect 45102 150618 64546 150854
rect 64782 150618 64866 150854
rect 65102 150618 84546 150854
rect 84782 150618 84866 150854
rect 85102 150618 104546 150854
rect 104782 150618 104866 150854
rect 105102 150618 124546 150854
rect 124782 150618 124866 150854
rect 125102 150618 144546 150854
rect 144782 150618 144866 150854
rect 145102 150618 164546 150854
rect 164782 150618 164866 150854
rect 165102 150618 184546 150854
rect 184782 150618 184866 150854
rect 185102 150618 204546 150854
rect 204782 150618 204866 150854
rect 205102 150618 224546 150854
rect 224782 150618 224866 150854
rect 225102 150618 244546 150854
rect 244782 150618 244866 150854
rect 245102 150618 264546 150854
rect 264782 150618 264866 150854
rect 265102 150618 284546 150854
rect 284782 150618 284866 150854
rect 285102 150618 304546 150854
rect 304782 150618 304866 150854
rect 305102 150618 324546 150854
rect 324782 150618 324866 150854
rect 325102 150618 344546 150854
rect 344782 150618 344866 150854
rect 345102 150618 364546 150854
rect 364782 150618 364866 150854
rect 365102 150618 384546 150854
rect 384782 150618 384866 150854
rect 385102 150618 404546 150854
rect 404782 150618 404866 150854
rect 405102 150618 424546 150854
rect 424782 150618 424866 150854
rect 425102 150618 444546 150854
rect 444782 150618 444866 150854
rect 445102 150618 464546 150854
rect 464782 150618 464866 150854
rect 465102 150618 484546 150854
rect 484782 150618 484866 150854
rect 485102 150618 504546 150854
rect 504782 150618 504866 150854
rect 505102 150618 524546 150854
rect 524782 150618 524866 150854
rect 525102 150618 544546 150854
rect 544782 150618 544866 150854
rect 545102 150618 564546 150854
rect 564782 150618 564866 150854
rect 565102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 826 147454
rect 1062 147218 1146 147454
rect 1382 147218 20826 147454
rect 21062 147218 21146 147454
rect 21382 147218 40826 147454
rect 41062 147218 41146 147454
rect 41382 147218 60826 147454
rect 61062 147218 61146 147454
rect 61382 147218 80826 147454
rect 81062 147218 81146 147454
rect 81382 147218 100826 147454
rect 101062 147218 101146 147454
rect 101382 147218 120826 147454
rect 121062 147218 121146 147454
rect 121382 147218 140826 147454
rect 141062 147218 141146 147454
rect 141382 147218 160826 147454
rect 161062 147218 161146 147454
rect 161382 147218 180826 147454
rect 181062 147218 181146 147454
rect 181382 147218 200826 147454
rect 201062 147218 201146 147454
rect 201382 147218 220826 147454
rect 221062 147218 221146 147454
rect 221382 147218 240826 147454
rect 241062 147218 241146 147454
rect 241382 147218 260826 147454
rect 261062 147218 261146 147454
rect 261382 147218 280826 147454
rect 281062 147218 281146 147454
rect 281382 147218 300826 147454
rect 301062 147218 301146 147454
rect 301382 147218 320826 147454
rect 321062 147218 321146 147454
rect 321382 147218 340826 147454
rect 341062 147218 341146 147454
rect 341382 147218 360826 147454
rect 361062 147218 361146 147454
rect 361382 147218 380826 147454
rect 381062 147218 381146 147454
rect 381382 147218 400826 147454
rect 401062 147218 401146 147454
rect 401382 147218 420826 147454
rect 421062 147218 421146 147454
rect 421382 147218 440826 147454
rect 441062 147218 441146 147454
rect 441382 147218 460826 147454
rect 461062 147218 461146 147454
rect 461382 147218 480826 147454
rect 481062 147218 481146 147454
rect 481382 147218 500826 147454
rect 501062 147218 501146 147454
rect 501382 147218 520826 147454
rect 521062 147218 521146 147454
rect 521382 147218 540826 147454
rect 541062 147218 541146 147454
rect 541382 147218 560826 147454
rect 561062 147218 561146 147454
rect 561382 147218 580826 147454
rect 581062 147218 581146 147454
rect 581382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 826 147134
rect 1062 146898 1146 147134
rect 1382 146898 20826 147134
rect 21062 146898 21146 147134
rect 21382 146898 40826 147134
rect 41062 146898 41146 147134
rect 41382 146898 60826 147134
rect 61062 146898 61146 147134
rect 61382 146898 80826 147134
rect 81062 146898 81146 147134
rect 81382 146898 100826 147134
rect 101062 146898 101146 147134
rect 101382 146898 120826 147134
rect 121062 146898 121146 147134
rect 121382 146898 140826 147134
rect 141062 146898 141146 147134
rect 141382 146898 160826 147134
rect 161062 146898 161146 147134
rect 161382 146898 180826 147134
rect 181062 146898 181146 147134
rect 181382 146898 200826 147134
rect 201062 146898 201146 147134
rect 201382 146898 220826 147134
rect 221062 146898 221146 147134
rect 221382 146898 240826 147134
rect 241062 146898 241146 147134
rect 241382 146898 260826 147134
rect 261062 146898 261146 147134
rect 261382 146898 280826 147134
rect 281062 146898 281146 147134
rect 281382 146898 300826 147134
rect 301062 146898 301146 147134
rect 301382 146898 320826 147134
rect 321062 146898 321146 147134
rect 321382 146898 340826 147134
rect 341062 146898 341146 147134
rect 341382 146898 360826 147134
rect 361062 146898 361146 147134
rect 361382 146898 380826 147134
rect 381062 146898 381146 147134
rect 381382 146898 400826 147134
rect 401062 146898 401146 147134
rect 401382 146898 420826 147134
rect 421062 146898 421146 147134
rect 421382 146898 440826 147134
rect 441062 146898 441146 147134
rect 441382 146898 460826 147134
rect 461062 146898 461146 147134
rect 461382 146898 480826 147134
rect 481062 146898 481146 147134
rect 481382 146898 500826 147134
rect 501062 146898 501146 147134
rect 501382 146898 520826 147134
rect 521062 146898 521146 147134
rect 521382 146898 540826 147134
rect 541062 146898 541146 147134
rect 541382 146898 560826 147134
rect 561062 146898 561146 147134
rect 561382 146898 580826 147134
rect 581062 146898 581146 147134
rect 581382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 21986 140614
rect 22222 140378 22306 140614
rect 22542 140378 41986 140614
rect 42222 140378 42306 140614
rect 42542 140378 61986 140614
rect 62222 140378 62306 140614
rect 62542 140378 81986 140614
rect 82222 140378 82306 140614
rect 82542 140378 101986 140614
rect 102222 140378 102306 140614
rect 102542 140378 121986 140614
rect 122222 140378 122306 140614
rect 122542 140378 141986 140614
rect 142222 140378 142306 140614
rect 142542 140378 161986 140614
rect 162222 140378 162306 140614
rect 162542 140378 181986 140614
rect 182222 140378 182306 140614
rect 182542 140378 201986 140614
rect 202222 140378 202306 140614
rect 202542 140378 221986 140614
rect 222222 140378 222306 140614
rect 222542 140378 241986 140614
rect 242222 140378 242306 140614
rect 242542 140378 261986 140614
rect 262222 140378 262306 140614
rect 262542 140378 281986 140614
rect 282222 140378 282306 140614
rect 282542 140378 301986 140614
rect 302222 140378 302306 140614
rect 302542 140378 321986 140614
rect 322222 140378 322306 140614
rect 322542 140378 341986 140614
rect 342222 140378 342306 140614
rect 342542 140378 361986 140614
rect 362222 140378 362306 140614
rect 362542 140378 381986 140614
rect 382222 140378 382306 140614
rect 382542 140378 401986 140614
rect 402222 140378 402306 140614
rect 402542 140378 421986 140614
rect 422222 140378 422306 140614
rect 422542 140378 441986 140614
rect 442222 140378 442306 140614
rect 442542 140378 461986 140614
rect 462222 140378 462306 140614
rect 462542 140378 481986 140614
rect 482222 140378 482306 140614
rect 482542 140378 501986 140614
rect 502222 140378 502306 140614
rect 502542 140378 521986 140614
rect 522222 140378 522306 140614
rect 522542 140378 541986 140614
rect 542222 140378 542306 140614
rect 542542 140378 561986 140614
rect 562222 140378 562306 140614
rect 562542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 21986 140294
rect 22222 140058 22306 140294
rect 22542 140058 41986 140294
rect 42222 140058 42306 140294
rect 42542 140058 61986 140294
rect 62222 140058 62306 140294
rect 62542 140058 81986 140294
rect 82222 140058 82306 140294
rect 82542 140058 101986 140294
rect 102222 140058 102306 140294
rect 102542 140058 121986 140294
rect 122222 140058 122306 140294
rect 122542 140058 141986 140294
rect 142222 140058 142306 140294
rect 142542 140058 161986 140294
rect 162222 140058 162306 140294
rect 162542 140058 181986 140294
rect 182222 140058 182306 140294
rect 182542 140058 201986 140294
rect 202222 140058 202306 140294
rect 202542 140058 221986 140294
rect 222222 140058 222306 140294
rect 222542 140058 241986 140294
rect 242222 140058 242306 140294
rect 242542 140058 261986 140294
rect 262222 140058 262306 140294
rect 262542 140058 281986 140294
rect 282222 140058 282306 140294
rect 282542 140058 301986 140294
rect 302222 140058 302306 140294
rect 302542 140058 321986 140294
rect 322222 140058 322306 140294
rect 322542 140058 341986 140294
rect 342222 140058 342306 140294
rect 342542 140058 361986 140294
rect 362222 140058 362306 140294
rect 362542 140058 381986 140294
rect 382222 140058 382306 140294
rect 382542 140058 401986 140294
rect 402222 140058 402306 140294
rect 402542 140058 421986 140294
rect 422222 140058 422306 140294
rect 422542 140058 441986 140294
rect 442222 140058 442306 140294
rect 442542 140058 461986 140294
rect 462222 140058 462306 140294
rect 462542 140058 481986 140294
rect 482222 140058 482306 140294
rect 482542 140058 501986 140294
rect 502222 140058 502306 140294
rect 502542 140058 521986 140294
rect 522222 140058 522306 140294
rect 522542 140058 541986 140294
rect 542222 140058 542306 140294
rect 542542 140058 561986 140294
rect 562222 140058 562306 140294
rect 562542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 18266 136894
rect 18502 136658 18586 136894
rect 18822 136658 38266 136894
rect 38502 136658 38586 136894
rect 38822 136658 58266 136894
rect 58502 136658 58586 136894
rect 58822 136658 78266 136894
rect 78502 136658 78586 136894
rect 78822 136658 98266 136894
rect 98502 136658 98586 136894
rect 98822 136658 118266 136894
rect 118502 136658 118586 136894
rect 118822 136658 138266 136894
rect 138502 136658 138586 136894
rect 138822 136658 158266 136894
rect 158502 136658 158586 136894
rect 158822 136658 178266 136894
rect 178502 136658 178586 136894
rect 178822 136658 198266 136894
rect 198502 136658 198586 136894
rect 198822 136658 218266 136894
rect 218502 136658 218586 136894
rect 218822 136658 238266 136894
rect 238502 136658 238586 136894
rect 238822 136658 258266 136894
rect 258502 136658 258586 136894
rect 258822 136658 278266 136894
rect 278502 136658 278586 136894
rect 278822 136658 298266 136894
rect 298502 136658 298586 136894
rect 298822 136658 318266 136894
rect 318502 136658 318586 136894
rect 318822 136658 338266 136894
rect 338502 136658 338586 136894
rect 338822 136658 358266 136894
rect 358502 136658 358586 136894
rect 358822 136658 378266 136894
rect 378502 136658 378586 136894
rect 378822 136658 398266 136894
rect 398502 136658 398586 136894
rect 398822 136658 418266 136894
rect 418502 136658 418586 136894
rect 418822 136658 438266 136894
rect 438502 136658 438586 136894
rect 438822 136658 458266 136894
rect 458502 136658 458586 136894
rect 458822 136658 478266 136894
rect 478502 136658 478586 136894
rect 478822 136658 498266 136894
rect 498502 136658 498586 136894
rect 498822 136658 518266 136894
rect 518502 136658 518586 136894
rect 518822 136658 538266 136894
rect 538502 136658 538586 136894
rect 538822 136658 558266 136894
rect 558502 136658 558586 136894
rect 558822 136658 578266 136894
rect 578502 136658 578586 136894
rect 578822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 18266 136574
rect 18502 136338 18586 136574
rect 18822 136338 38266 136574
rect 38502 136338 38586 136574
rect 38822 136338 58266 136574
rect 58502 136338 58586 136574
rect 58822 136338 78266 136574
rect 78502 136338 78586 136574
rect 78822 136338 98266 136574
rect 98502 136338 98586 136574
rect 98822 136338 118266 136574
rect 118502 136338 118586 136574
rect 118822 136338 138266 136574
rect 138502 136338 138586 136574
rect 138822 136338 158266 136574
rect 158502 136338 158586 136574
rect 158822 136338 178266 136574
rect 178502 136338 178586 136574
rect 178822 136338 198266 136574
rect 198502 136338 198586 136574
rect 198822 136338 218266 136574
rect 218502 136338 218586 136574
rect 218822 136338 238266 136574
rect 238502 136338 238586 136574
rect 238822 136338 258266 136574
rect 258502 136338 258586 136574
rect 258822 136338 278266 136574
rect 278502 136338 278586 136574
rect 278822 136338 298266 136574
rect 298502 136338 298586 136574
rect 298822 136338 318266 136574
rect 318502 136338 318586 136574
rect 318822 136338 338266 136574
rect 338502 136338 338586 136574
rect 338822 136338 358266 136574
rect 358502 136338 358586 136574
rect 358822 136338 378266 136574
rect 378502 136338 378586 136574
rect 378822 136338 398266 136574
rect 398502 136338 398586 136574
rect 398822 136338 418266 136574
rect 418502 136338 418586 136574
rect 418822 136338 438266 136574
rect 438502 136338 438586 136574
rect 438822 136338 458266 136574
rect 458502 136338 458586 136574
rect 458822 136338 478266 136574
rect 478502 136338 478586 136574
rect 478822 136338 498266 136574
rect 498502 136338 498586 136574
rect 498822 136338 518266 136574
rect 518502 136338 518586 136574
rect 518822 136338 538266 136574
rect 538502 136338 538586 136574
rect 538822 136338 558266 136574
rect 558502 136338 558586 136574
rect 558822 136338 578266 136574
rect 578502 136338 578586 136574
rect 578822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 14546 133174
rect 14782 132938 14866 133174
rect 15102 132938 34546 133174
rect 34782 132938 34866 133174
rect 35102 132938 54546 133174
rect 54782 132938 54866 133174
rect 55102 132938 74546 133174
rect 74782 132938 74866 133174
rect 75102 132938 94546 133174
rect 94782 132938 94866 133174
rect 95102 132938 114546 133174
rect 114782 132938 114866 133174
rect 115102 132938 134546 133174
rect 134782 132938 134866 133174
rect 135102 132938 154546 133174
rect 154782 132938 154866 133174
rect 155102 132938 174546 133174
rect 174782 132938 174866 133174
rect 175102 132938 194546 133174
rect 194782 132938 194866 133174
rect 195102 132938 214546 133174
rect 214782 132938 214866 133174
rect 215102 132938 234546 133174
rect 234782 132938 234866 133174
rect 235102 132938 254546 133174
rect 254782 132938 254866 133174
rect 255102 132938 274546 133174
rect 274782 132938 274866 133174
rect 275102 132938 294546 133174
rect 294782 132938 294866 133174
rect 295102 132938 314546 133174
rect 314782 132938 314866 133174
rect 315102 132938 334546 133174
rect 334782 132938 334866 133174
rect 335102 132938 354546 133174
rect 354782 132938 354866 133174
rect 355102 132938 374546 133174
rect 374782 132938 374866 133174
rect 375102 132938 394546 133174
rect 394782 132938 394866 133174
rect 395102 132938 414546 133174
rect 414782 132938 414866 133174
rect 415102 132938 434546 133174
rect 434782 132938 434866 133174
rect 435102 132938 454546 133174
rect 454782 132938 454866 133174
rect 455102 132938 474546 133174
rect 474782 132938 474866 133174
rect 475102 132938 494546 133174
rect 494782 132938 494866 133174
rect 495102 132938 514546 133174
rect 514782 132938 514866 133174
rect 515102 132938 534546 133174
rect 534782 132938 534866 133174
rect 535102 132938 554546 133174
rect 554782 132938 554866 133174
rect 555102 132938 574546 133174
rect 574782 132938 574866 133174
rect 575102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 14546 132854
rect 14782 132618 14866 132854
rect 15102 132618 34546 132854
rect 34782 132618 34866 132854
rect 35102 132618 54546 132854
rect 54782 132618 54866 132854
rect 55102 132618 74546 132854
rect 74782 132618 74866 132854
rect 75102 132618 94546 132854
rect 94782 132618 94866 132854
rect 95102 132618 114546 132854
rect 114782 132618 114866 132854
rect 115102 132618 134546 132854
rect 134782 132618 134866 132854
rect 135102 132618 154546 132854
rect 154782 132618 154866 132854
rect 155102 132618 174546 132854
rect 174782 132618 174866 132854
rect 175102 132618 194546 132854
rect 194782 132618 194866 132854
rect 195102 132618 214546 132854
rect 214782 132618 214866 132854
rect 215102 132618 234546 132854
rect 234782 132618 234866 132854
rect 235102 132618 254546 132854
rect 254782 132618 254866 132854
rect 255102 132618 274546 132854
rect 274782 132618 274866 132854
rect 275102 132618 294546 132854
rect 294782 132618 294866 132854
rect 295102 132618 314546 132854
rect 314782 132618 314866 132854
rect 315102 132618 334546 132854
rect 334782 132618 334866 132854
rect 335102 132618 354546 132854
rect 354782 132618 354866 132854
rect 355102 132618 374546 132854
rect 374782 132618 374866 132854
rect 375102 132618 394546 132854
rect 394782 132618 394866 132854
rect 395102 132618 414546 132854
rect 414782 132618 414866 132854
rect 415102 132618 434546 132854
rect 434782 132618 434866 132854
rect 435102 132618 454546 132854
rect 454782 132618 454866 132854
rect 455102 132618 474546 132854
rect 474782 132618 474866 132854
rect 475102 132618 494546 132854
rect 494782 132618 494866 132854
rect 495102 132618 514546 132854
rect 514782 132618 514866 132854
rect 515102 132618 534546 132854
rect 534782 132618 534866 132854
rect 535102 132618 554546 132854
rect 554782 132618 554866 132854
rect 555102 132618 574546 132854
rect 574782 132618 574866 132854
rect 575102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 10826 129454
rect 11062 129218 11146 129454
rect 11382 129218 30826 129454
rect 31062 129218 31146 129454
rect 31382 129218 50826 129454
rect 51062 129218 51146 129454
rect 51382 129218 70826 129454
rect 71062 129218 71146 129454
rect 71382 129218 90826 129454
rect 91062 129218 91146 129454
rect 91382 129218 110826 129454
rect 111062 129218 111146 129454
rect 111382 129218 130826 129454
rect 131062 129218 131146 129454
rect 131382 129218 150826 129454
rect 151062 129218 151146 129454
rect 151382 129218 170826 129454
rect 171062 129218 171146 129454
rect 171382 129218 190826 129454
rect 191062 129218 191146 129454
rect 191382 129218 210826 129454
rect 211062 129218 211146 129454
rect 211382 129218 230826 129454
rect 231062 129218 231146 129454
rect 231382 129218 250826 129454
rect 251062 129218 251146 129454
rect 251382 129218 270826 129454
rect 271062 129218 271146 129454
rect 271382 129218 290826 129454
rect 291062 129218 291146 129454
rect 291382 129218 310826 129454
rect 311062 129218 311146 129454
rect 311382 129218 330826 129454
rect 331062 129218 331146 129454
rect 331382 129218 350826 129454
rect 351062 129218 351146 129454
rect 351382 129218 370826 129454
rect 371062 129218 371146 129454
rect 371382 129218 390826 129454
rect 391062 129218 391146 129454
rect 391382 129218 410826 129454
rect 411062 129218 411146 129454
rect 411382 129218 430826 129454
rect 431062 129218 431146 129454
rect 431382 129218 450826 129454
rect 451062 129218 451146 129454
rect 451382 129218 470826 129454
rect 471062 129218 471146 129454
rect 471382 129218 490826 129454
rect 491062 129218 491146 129454
rect 491382 129218 510826 129454
rect 511062 129218 511146 129454
rect 511382 129218 530826 129454
rect 531062 129218 531146 129454
rect 531382 129218 550826 129454
rect 551062 129218 551146 129454
rect 551382 129218 570826 129454
rect 571062 129218 571146 129454
rect 571382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 10826 129134
rect 11062 128898 11146 129134
rect 11382 128898 30826 129134
rect 31062 128898 31146 129134
rect 31382 128898 50826 129134
rect 51062 128898 51146 129134
rect 51382 128898 70826 129134
rect 71062 128898 71146 129134
rect 71382 128898 90826 129134
rect 91062 128898 91146 129134
rect 91382 128898 110826 129134
rect 111062 128898 111146 129134
rect 111382 128898 130826 129134
rect 131062 128898 131146 129134
rect 131382 128898 150826 129134
rect 151062 128898 151146 129134
rect 151382 128898 170826 129134
rect 171062 128898 171146 129134
rect 171382 128898 190826 129134
rect 191062 128898 191146 129134
rect 191382 128898 210826 129134
rect 211062 128898 211146 129134
rect 211382 128898 230826 129134
rect 231062 128898 231146 129134
rect 231382 128898 250826 129134
rect 251062 128898 251146 129134
rect 251382 128898 270826 129134
rect 271062 128898 271146 129134
rect 271382 128898 290826 129134
rect 291062 128898 291146 129134
rect 291382 128898 310826 129134
rect 311062 128898 311146 129134
rect 311382 128898 330826 129134
rect 331062 128898 331146 129134
rect 331382 128898 350826 129134
rect 351062 128898 351146 129134
rect 351382 128898 370826 129134
rect 371062 128898 371146 129134
rect 371382 128898 390826 129134
rect 391062 128898 391146 129134
rect 391382 128898 410826 129134
rect 411062 128898 411146 129134
rect 411382 128898 430826 129134
rect 431062 128898 431146 129134
rect 431382 128898 450826 129134
rect 451062 128898 451146 129134
rect 451382 128898 470826 129134
rect 471062 128898 471146 129134
rect 471382 128898 490826 129134
rect 491062 128898 491146 129134
rect 491382 128898 510826 129134
rect 511062 128898 511146 129134
rect 511382 128898 530826 129134
rect 531062 128898 531146 129134
rect 531382 128898 550826 129134
rect 551062 128898 551146 129134
rect 551382 128898 570826 129134
rect 571062 128898 571146 129134
rect 571382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 11986 122614
rect 12222 122378 12306 122614
rect 12542 122378 31986 122614
rect 32222 122378 32306 122614
rect 32542 122378 51986 122614
rect 52222 122378 52306 122614
rect 52542 122378 71986 122614
rect 72222 122378 72306 122614
rect 72542 122378 91986 122614
rect 92222 122378 92306 122614
rect 92542 122378 111986 122614
rect 112222 122378 112306 122614
rect 112542 122378 131986 122614
rect 132222 122378 132306 122614
rect 132542 122378 151986 122614
rect 152222 122378 152306 122614
rect 152542 122378 171986 122614
rect 172222 122378 172306 122614
rect 172542 122378 191986 122614
rect 192222 122378 192306 122614
rect 192542 122378 211986 122614
rect 212222 122378 212306 122614
rect 212542 122378 231986 122614
rect 232222 122378 232306 122614
rect 232542 122378 251986 122614
rect 252222 122378 252306 122614
rect 252542 122378 271986 122614
rect 272222 122378 272306 122614
rect 272542 122378 291986 122614
rect 292222 122378 292306 122614
rect 292542 122378 311986 122614
rect 312222 122378 312306 122614
rect 312542 122378 331986 122614
rect 332222 122378 332306 122614
rect 332542 122378 351986 122614
rect 352222 122378 352306 122614
rect 352542 122378 371986 122614
rect 372222 122378 372306 122614
rect 372542 122378 391986 122614
rect 392222 122378 392306 122614
rect 392542 122378 411986 122614
rect 412222 122378 412306 122614
rect 412542 122378 431986 122614
rect 432222 122378 432306 122614
rect 432542 122378 451986 122614
rect 452222 122378 452306 122614
rect 452542 122378 471986 122614
rect 472222 122378 472306 122614
rect 472542 122378 491986 122614
rect 492222 122378 492306 122614
rect 492542 122378 511986 122614
rect 512222 122378 512306 122614
rect 512542 122378 531986 122614
rect 532222 122378 532306 122614
rect 532542 122378 551986 122614
rect 552222 122378 552306 122614
rect 552542 122378 571986 122614
rect 572222 122378 572306 122614
rect 572542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 11986 122294
rect 12222 122058 12306 122294
rect 12542 122058 31986 122294
rect 32222 122058 32306 122294
rect 32542 122058 51986 122294
rect 52222 122058 52306 122294
rect 52542 122058 71986 122294
rect 72222 122058 72306 122294
rect 72542 122058 91986 122294
rect 92222 122058 92306 122294
rect 92542 122058 111986 122294
rect 112222 122058 112306 122294
rect 112542 122058 131986 122294
rect 132222 122058 132306 122294
rect 132542 122058 151986 122294
rect 152222 122058 152306 122294
rect 152542 122058 171986 122294
rect 172222 122058 172306 122294
rect 172542 122058 191986 122294
rect 192222 122058 192306 122294
rect 192542 122058 211986 122294
rect 212222 122058 212306 122294
rect 212542 122058 231986 122294
rect 232222 122058 232306 122294
rect 232542 122058 251986 122294
rect 252222 122058 252306 122294
rect 252542 122058 271986 122294
rect 272222 122058 272306 122294
rect 272542 122058 291986 122294
rect 292222 122058 292306 122294
rect 292542 122058 311986 122294
rect 312222 122058 312306 122294
rect 312542 122058 331986 122294
rect 332222 122058 332306 122294
rect 332542 122058 351986 122294
rect 352222 122058 352306 122294
rect 352542 122058 371986 122294
rect 372222 122058 372306 122294
rect 372542 122058 391986 122294
rect 392222 122058 392306 122294
rect 392542 122058 411986 122294
rect 412222 122058 412306 122294
rect 412542 122058 431986 122294
rect 432222 122058 432306 122294
rect 432542 122058 451986 122294
rect 452222 122058 452306 122294
rect 452542 122058 471986 122294
rect 472222 122058 472306 122294
rect 472542 122058 491986 122294
rect 492222 122058 492306 122294
rect 492542 122058 511986 122294
rect 512222 122058 512306 122294
rect 512542 122058 531986 122294
rect 532222 122058 532306 122294
rect 532542 122058 551986 122294
rect 552222 122058 552306 122294
rect 552542 122058 571986 122294
rect 572222 122058 572306 122294
rect 572542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 8266 118894
rect 8502 118658 8586 118894
rect 8822 118658 28266 118894
rect 28502 118658 28586 118894
rect 28822 118658 48266 118894
rect 48502 118658 48586 118894
rect 48822 118658 68266 118894
rect 68502 118658 68586 118894
rect 68822 118658 88266 118894
rect 88502 118658 88586 118894
rect 88822 118658 108266 118894
rect 108502 118658 108586 118894
rect 108822 118658 128266 118894
rect 128502 118658 128586 118894
rect 128822 118658 148266 118894
rect 148502 118658 148586 118894
rect 148822 118658 168266 118894
rect 168502 118658 168586 118894
rect 168822 118658 188266 118894
rect 188502 118658 188586 118894
rect 188822 118658 208266 118894
rect 208502 118658 208586 118894
rect 208822 118658 228266 118894
rect 228502 118658 228586 118894
rect 228822 118658 248266 118894
rect 248502 118658 248586 118894
rect 248822 118658 268266 118894
rect 268502 118658 268586 118894
rect 268822 118658 288266 118894
rect 288502 118658 288586 118894
rect 288822 118658 308266 118894
rect 308502 118658 308586 118894
rect 308822 118658 328266 118894
rect 328502 118658 328586 118894
rect 328822 118658 348266 118894
rect 348502 118658 348586 118894
rect 348822 118658 368266 118894
rect 368502 118658 368586 118894
rect 368822 118658 388266 118894
rect 388502 118658 388586 118894
rect 388822 118658 408266 118894
rect 408502 118658 408586 118894
rect 408822 118658 428266 118894
rect 428502 118658 428586 118894
rect 428822 118658 448266 118894
rect 448502 118658 448586 118894
rect 448822 118658 468266 118894
rect 468502 118658 468586 118894
rect 468822 118658 488266 118894
rect 488502 118658 488586 118894
rect 488822 118658 508266 118894
rect 508502 118658 508586 118894
rect 508822 118658 528266 118894
rect 528502 118658 528586 118894
rect 528822 118658 548266 118894
rect 548502 118658 548586 118894
rect 548822 118658 568266 118894
rect 568502 118658 568586 118894
rect 568822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 8266 118574
rect 8502 118338 8586 118574
rect 8822 118338 28266 118574
rect 28502 118338 28586 118574
rect 28822 118338 48266 118574
rect 48502 118338 48586 118574
rect 48822 118338 68266 118574
rect 68502 118338 68586 118574
rect 68822 118338 88266 118574
rect 88502 118338 88586 118574
rect 88822 118338 108266 118574
rect 108502 118338 108586 118574
rect 108822 118338 128266 118574
rect 128502 118338 128586 118574
rect 128822 118338 148266 118574
rect 148502 118338 148586 118574
rect 148822 118338 168266 118574
rect 168502 118338 168586 118574
rect 168822 118338 188266 118574
rect 188502 118338 188586 118574
rect 188822 118338 208266 118574
rect 208502 118338 208586 118574
rect 208822 118338 228266 118574
rect 228502 118338 228586 118574
rect 228822 118338 248266 118574
rect 248502 118338 248586 118574
rect 248822 118338 268266 118574
rect 268502 118338 268586 118574
rect 268822 118338 288266 118574
rect 288502 118338 288586 118574
rect 288822 118338 308266 118574
rect 308502 118338 308586 118574
rect 308822 118338 328266 118574
rect 328502 118338 328586 118574
rect 328822 118338 348266 118574
rect 348502 118338 348586 118574
rect 348822 118338 368266 118574
rect 368502 118338 368586 118574
rect 368822 118338 388266 118574
rect 388502 118338 388586 118574
rect 388822 118338 408266 118574
rect 408502 118338 408586 118574
rect 408822 118338 428266 118574
rect 428502 118338 428586 118574
rect 428822 118338 448266 118574
rect 448502 118338 448586 118574
rect 448822 118338 468266 118574
rect 468502 118338 468586 118574
rect 468822 118338 488266 118574
rect 488502 118338 488586 118574
rect 488822 118338 508266 118574
rect 508502 118338 508586 118574
rect 508822 118338 528266 118574
rect 528502 118338 528586 118574
rect 528822 118338 548266 118574
rect 548502 118338 548586 118574
rect 548822 118338 568266 118574
rect 568502 118338 568586 118574
rect 568822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 4546 115174
rect 4782 114938 4866 115174
rect 5102 114938 24546 115174
rect 24782 114938 24866 115174
rect 25102 114938 44546 115174
rect 44782 114938 44866 115174
rect 45102 114938 64546 115174
rect 64782 114938 64866 115174
rect 65102 114938 84546 115174
rect 84782 114938 84866 115174
rect 85102 114938 104546 115174
rect 104782 114938 104866 115174
rect 105102 114938 124546 115174
rect 124782 114938 124866 115174
rect 125102 114938 144546 115174
rect 144782 114938 144866 115174
rect 145102 114938 164546 115174
rect 164782 114938 164866 115174
rect 165102 114938 184546 115174
rect 184782 114938 184866 115174
rect 185102 114938 204546 115174
rect 204782 114938 204866 115174
rect 205102 114938 224546 115174
rect 224782 114938 224866 115174
rect 225102 114938 244546 115174
rect 244782 114938 244866 115174
rect 245102 114938 264546 115174
rect 264782 114938 264866 115174
rect 265102 114938 284546 115174
rect 284782 114938 284866 115174
rect 285102 114938 304546 115174
rect 304782 114938 304866 115174
rect 305102 114938 324546 115174
rect 324782 114938 324866 115174
rect 325102 114938 344546 115174
rect 344782 114938 344866 115174
rect 345102 114938 364546 115174
rect 364782 114938 364866 115174
rect 365102 114938 384546 115174
rect 384782 114938 384866 115174
rect 385102 114938 404546 115174
rect 404782 114938 404866 115174
rect 405102 114938 424546 115174
rect 424782 114938 424866 115174
rect 425102 114938 444546 115174
rect 444782 114938 444866 115174
rect 445102 114938 464546 115174
rect 464782 114938 464866 115174
rect 465102 114938 484546 115174
rect 484782 114938 484866 115174
rect 485102 114938 504546 115174
rect 504782 114938 504866 115174
rect 505102 114938 524546 115174
rect 524782 114938 524866 115174
rect 525102 114938 544546 115174
rect 544782 114938 544866 115174
rect 545102 114938 564546 115174
rect 564782 114938 564866 115174
rect 565102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 4546 114854
rect 4782 114618 4866 114854
rect 5102 114618 24546 114854
rect 24782 114618 24866 114854
rect 25102 114618 44546 114854
rect 44782 114618 44866 114854
rect 45102 114618 64546 114854
rect 64782 114618 64866 114854
rect 65102 114618 84546 114854
rect 84782 114618 84866 114854
rect 85102 114618 104546 114854
rect 104782 114618 104866 114854
rect 105102 114618 124546 114854
rect 124782 114618 124866 114854
rect 125102 114618 144546 114854
rect 144782 114618 144866 114854
rect 145102 114618 164546 114854
rect 164782 114618 164866 114854
rect 165102 114618 184546 114854
rect 184782 114618 184866 114854
rect 185102 114618 204546 114854
rect 204782 114618 204866 114854
rect 205102 114618 224546 114854
rect 224782 114618 224866 114854
rect 225102 114618 244546 114854
rect 244782 114618 244866 114854
rect 245102 114618 264546 114854
rect 264782 114618 264866 114854
rect 265102 114618 284546 114854
rect 284782 114618 284866 114854
rect 285102 114618 304546 114854
rect 304782 114618 304866 114854
rect 305102 114618 324546 114854
rect 324782 114618 324866 114854
rect 325102 114618 344546 114854
rect 344782 114618 344866 114854
rect 345102 114618 364546 114854
rect 364782 114618 364866 114854
rect 365102 114618 384546 114854
rect 384782 114618 384866 114854
rect 385102 114618 404546 114854
rect 404782 114618 404866 114854
rect 405102 114618 424546 114854
rect 424782 114618 424866 114854
rect 425102 114618 444546 114854
rect 444782 114618 444866 114854
rect 445102 114618 464546 114854
rect 464782 114618 464866 114854
rect 465102 114618 484546 114854
rect 484782 114618 484866 114854
rect 485102 114618 504546 114854
rect 504782 114618 504866 114854
rect 505102 114618 524546 114854
rect 524782 114618 524866 114854
rect 525102 114618 544546 114854
rect 544782 114618 544866 114854
rect 545102 114618 564546 114854
rect 564782 114618 564866 114854
rect 565102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 826 111454
rect 1062 111218 1146 111454
rect 1382 111218 20826 111454
rect 21062 111218 21146 111454
rect 21382 111218 40826 111454
rect 41062 111218 41146 111454
rect 41382 111218 60826 111454
rect 61062 111218 61146 111454
rect 61382 111218 80826 111454
rect 81062 111218 81146 111454
rect 81382 111218 100826 111454
rect 101062 111218 101146 111454
rect 101382 111218 120826 111454
rect 121062 111218 121146 111454
rect 121382 111218 140826 111454
rect 141062 111218 141146 111454
rect 141382 111218 160826 111454
rect 161062 111218 161146 111454
rect 161382 111218 180826 111454
rect 181062 111218 181146 111454
rect 181382 111218 200826 111454
rect 201062 111218 201146 111454
rect 201382 111218 220826 111454
rect 221062 111218 221146 111454
rect 221382 111218 240826 111454
rect 241062 111218 241146 111454
rect 241382 111218 260826 111454
rect 261062 111218 261146 111454
rect 261382 111218 280826 111454
rect 281062 111218 281146 111454
rect 281382 111218 300826 111454
rect 301062 111218 301146 111454
rect 301382 111218 320826 111454
rect 321062 111218 321146 111454
rect 321382 111218 340826 111454
rect 341062 111218 341146 111454
rect 341382 111218 360826 111454
rect 361062 111218 361146 111454
rect 361382 111218 380826 111454
rect 381062 111218 381146 111454
rect 381382 111218 400826 111454
rect 401062 111218 401146 111454
rect 401382 111218 420826 111454
rect 421062 111218 421146 111454
rect 421382 111218 440826 111454
rect 441062 111218 441146 111454
rect 441382 111218 460826 111454
rect 461062 111218 461146 111454
rect 461382 111218 480826 111454
rect 481062 111218 481146 111454
rect 481382 111218 500826 111454
rect 501062 111218 501146 111454
rect 501382 111218 520826 111454
rect 521062 111218 521146 111454
rect 521382 111218 540826 111454
rect 541062 111218 541146 111454
rect 541382 111218 560826 111454
rect 561062 111218 561146 111454
rect 561382 111218 580826 111454
rect 581062 111218 581146 111454
rect 581382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 826 111134
rect 1062 110898 1146 111134
rect 1382 110898 20826 111134
rect 21062 110898 21146 111134
rect 21382 110898 40826 111134
rect 41062 110898 41146 111134
rect 41382 110898 60826 111134
rect 61062 110898 61146 111134
rect 61382 110898 80826 111134
rect 81062 110898 81146 111134
rect 81382 110898 100826 111134
rect 101062 110898 101146 111134
rect 101382 110898 120826 111134
rect 121062 110898 121146 111134
rect 121382 110898 140826 111134
rect 141062 110898 141146 111134
rect 141382 110898 160826 111134
rect 161062 110898 161146 111134
rect 161382 110898 180826 111134
rect 181062 110898 181146 111134
rect 181382 110898 200826 111134
rect 201062 110898 201146 111134
rect 201382 110898 220826 111134
rect 221062 110898 221146 111134
rect 221382 110898 240826 111134
rect 241062 110898 241146 111134
rect 241382 110898 260826 111134
rect 261062 110898 261146 111134
rect 261382 110898 280826 111134
rect 281062 110898 281146 111134
rect 281382 110898 300826 111134
rect 301062 110898 301146 111134
rect 301382 110898 320826 111134
rect 321062 110898 321146 111134
rect 321382 110898 340826 111134
rect 341062 110898 341146 111134
rect 341382 110898 360826 111134
rect 361062 110898 361146 111134
rect 361382 110898 380826 111134
rect 381062 110898 381146 111134
rect 381382 110898 400826 111134
rect 401062 110898 401146 111134
rect 401382 110898 420826 111134
rect 421062 110898 421146 111134
rect 421382 110898 440826 111134
rect 441062 110898 441146 111134
rect 441382 110898 460826 111134
rect 461062 110898 461146 111134
rect 461382 110898 480826 111134
rect 481062 110898 481146 111134
rect 481382 110898 500826 111134
rect 501062 110898 501146 111134
rect 501382 110898 520826 111134
rect 521062 110898 521146 111134
rect 521382 110898 540826 111134
rect 541062 110898 541146 111134
rect 541382 110898 560826 111134
rect 561062 110898 561146 111134
rect 561382 110898 580826 111134
rect 581062 110898 581146 111134
rect 581382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 21986 104614
rect 22222 104378 22306 104614
rect 22542 104378 41986 104614
rect 42222 104378 42306 104614
rect 42542 104378 61986 104614
rect 62222 104378 62306 104614
rect 62542 104378 81986 104614
rect 82222 104378 82306 104614
rect 82542 104378 101986 104614
rect 102222 104378 102306 104614
rect 102542 104378 121986 104614
rect 122222 104378 122306 104614
rect 122542 104378 141986 104614
rect 142222 104378 142306 104614
rect 142542 104378 161986 104614
rect 162222 104378 162306 104614
rect 162542 104378 181986 104614
rect 182222 104378 182306 104614
rect 182542 104378 201986 104614
rect 202222 104378 202306 104614
rect 202542 104378 221986 104614
rect 222222 104378 222306 104614
rect 222542 104378 241986 104614
rect 242222 104378 242306 104614
rect 242542 104378 261986 104614
rect 262222 104378 262306 104614
rect 262542 104378 281986 104614
rect 282222 104378 282306 104614
rect 282542 104378 301986 104614
rect 302222 104378 302306 104614
rect 302542 104378 321986 104614
rect 322222 104378 322306 104614
rect 322542 104378 341986 104614
rect 342222 104378 342306 104614
rect 342542 104378 361986 104614
rect 362222 104378 362306 104614
rect 362542 104378 381986 104614
rect 382222 104378 382306 104614
rect 382542 104378 401986 104614
rect 402222 104378 402306 104614
rect 402542 104378 421986 104614
rect 422222 104378 422306 104614
rect 422542 104378 441986 104614
rect 442222 104378 442306 104614
rect 442542 104378 461986 104614
rect 462222 104378 462306 104614
rect 462542 104378 481986 104614
rect 482222 104378 482306 104614
rect 482542 104378 501986 104614
rect 502222 104378 502306 104614
rect 502542 104378 521986 104614
rect 522222 104378 522306 104614
rect 522542 104378 541986 104614
rect 542222 104378 542306 104614
rect 542542 104378 561986 104614
rect 562222 104378 562306 104614
rect 562542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 21986 104294
rect 22222 104058 22306 104294
rect 22542 104058 41986 104294
rect 42222 104058 42306 104294
rect 42542 104058 61986 104294
rect 62222 104058 62306 104294
rect 62542 104058 81986 104294
rect 82222 104058 82306 104294
rect 82542 104058 101986 104294
rect 102222 104058 102306 104294
rect 102542 104058 121986 104294
rect 122222 104058 122306 104294
rect 122542 104058 141986 104294
rect 142222 104058 142306 104294
rect 142542 104058 161986 104294
rect 162222 104058 162306 104294
rect 162542 104058 181986 104294
rect 182222 104058 182306 104294
rect 182542 104058 201986 104294
rect 202222 104058 202306 104294
rect 202542 104058 221986 104294
rect 222222 104058 222306 104294
rect 222542 104058 241986 104294
rect 242222 104058 242306 104294
rect 242542 104058 261986 104294
rect 262222 104058 262306 104294
rect 262542 104058 281986 104294
rect 282222 104058 282306 104294
rect 282542 104058 301986 104294
rect 302222 104058 302306 104294
rect 302542 104058 321986 104294
rect 322222 104058 322306 104294
rect 322542 104058 341986 104294
rect 342222 104058 342306 104294
rect 342542 104058 361986 104294
rect 362222 104058 362306 104294
rect 362542 104058 381986 104294
rect 382222 104058 382306 104294
rect 382542 104058 401986 104294
rect 402222 104058 402306 104294
rect 402542 104058 421986 104294
rect 422222 104058 422306 104294
rect 422542 104058 441986 104294
rect 442222 104058 442306 104294
rect 442542 104058 461986 104294
rect 462222 104058 462306 104294
rect 462542 104058 481986 104294
rect 482222 104058 482306 104294
rect 482542 104058 501986 104294
rect 502222 104058 502306 104294
rect 502542 104058 521986 104294
rect 522222 104058 522306 104294
rect 522542 104058 541986 104294
rect 542222 104058 542306 104294
rect 542542 104058 561986 104294
rect 562222 104058 562306 104294
rect 562542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 18266 100894
rect 18502 100658 18586 100894
rect 18822 100658 38266 100894
rect 38502 100658 38586 100894
rect 38822 100658 58266 100894
rect 58502 100658 58586 100894
rect 58822 100658 78266 100894
rect 78502 100658 78586 100894
rect 78822 100658 98266 100894
rect 98502 100658 98586 100894
rect 98822 100658 118266 100894
rect 118502 100658 118586 100894
rect 118822 100658 138266 100894
rect 138502 100658 138586 100894
rect 138822 100658 158266 100894
rect 158502 100658 158586 100894
rect 158822 100658 178266 100894
rect 178502 100658 178586 100894
rect 178822 100658 198266 100894
rect 198502 100658 198586 100894
rect 198822 100658 218266 100894
rect 218502 100658 218586 100894
rect 218822 100658 238266 100894
rect 238502 100658 238586 100894
rect 238822 100658 258266 100894
rect 258502 100658 258586 100894
rect 258822 100658 278266 100894
rect 278502 100658 278586 100894
rect 278822 100658 298266 100894
rect 298502 100658 298586 100894
rect 298822 100658 318266 100894
rect 318502 100658 318586 100894
rect 318822 100658 338266 100894
rect 338502 100658 338586 100894
rect 338822 100658 358266 100894
rect 358502 100658 358586 100894
rect 358822 100658 378266 100894
rect 378502 100658 378586 100894
rect 378822 100658 398266 100894
rect 398502 100658 398586 100894
rect 398822 100658 418266 100894
rect 418502 100658 418586 100894
rect 418822 100658 438266 100894
rect 438502 100658 438586 100894
rect 438822 100658 458266 100894
rect 458502 100658 458586 100894
rect 458822 100658 478266 100894
rect 478502 100658 478586 100894
rect 478822 100658 498266 100894
rect 498502 100658 498586 100894
rect 498822 100658 518266 100894
rect 518502 100658 518586 100894
rect 518822 100658 538266 100894
rect 538502 100658 538586 100894
rect 538822 100658 558266 100894
rect 558502 100658 558586 100894
rect 558822 100658 578266 100894
rect 578502 100658 578586 100894
rect 578822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 18266 100574
rect 18502 100338 18586 100574
rect 18822 100338 38266 100574
rect 38502 100338 38586 100574
rect 38822 100338 58266 100574
rect 58502 100338 58586 100574
rect 58822 100338 78266 100574
rect 78502 100338 78586 100574
rect 78822 100338 98266 100574
rect 98502 100338 98586 100574
rect 98822 100338 118266 100574
rect 118502 100338 118586 100574
rect 118822 100338 138266 100574
rect 138502 100338 138586 100574
rect 138822 100338 158266 100574
rect 158502 100338 158586 100574
rect 158822 100338 178266 100574
rect 178502 100338 178586 100574
rect 178822 100338 198266 100574
rect 198502 100338 198586 100574
rect 198822 100338 218266 100574
rect 218502 100338 218586 100574
rect 218822 100338 238266 100574
rect 238502 100338 238586 100574
rect 238822 100338 258266 100574
rect 258502 100338 258586 100574
rect 258822 100338 278266 100574
rect 278502 100338 278586 100574
rect 278822 100338 298266 100574
rect 298502 100338 298586 100574
rect 298822 100338 318266 100574
rect 318502 100338 318586 100574
rect 318822 100338 338266 100574
rect 338502 100338 338586 100574
rect 338822 100338 358266 100574
rect 358502 100338 358586 100574
rect 358822 100338 378266 100574
rect 378502 100338 378586 100574
rect 378822 100338 398266 100574
rect 398502 100338 398586 100574
rect 398822 100338 418266 100574
rect 418502 100338 418586 100574
rect 418822 100338 438266 100574
rect 438502 100338 438586 100574
rect 438822 100338 458266 100574
rect 458502 100338 458586 100574
rect 458822 100338 478266 100574
rect 478502 100338 478586 100574
rect 478822 100338 498266 100574
rect 498502 100338 498586 100574
rect 498822 100338 518266 100574
rect 518502 100338 518586 100574
rect 518822 100338 538266 100574
rect 538502 100338 538586 100574
rect 538822 100338 558266 100574
rect 558502 100338 558586 100574
rect 558822 100338 578266 100574
rect 578502 100338 578586 100574
rect 578822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 14546 97174
rect 14782 96938 14866 97174
rect 15102 96938 34546 97174
rect 34782 96938 34866 97174
rect 35102 96938 54546 97174
rect 54782 96938 54866 97174
rect 55102 96938 74546 97174
rect 74782 96938 74866 97174
rect 75102 96938 94546 97174
rect 94782 96938 94866 97174
rect 95102 96938 114546 97174
rect 114782 96938 114866 97174
rect 115102 96938 134546 97174
rect 134782 96938 134866 97174
rect 135102 96938 154546 97174
rect 154782 96938 154866 97174
rect 155102 96938 174546 97174
rect 174782 96938 174866 97174
rect 175102 96938 194546 97174
rect 194782 96938 194866 97174
rect 195102 96938 214546 97174
rect 214782 96938 214866 97174
rect 215102 96938 234546 97174
rect 234782 96938 234866 97174
rect 235102 96938 254546 97174
rect 254782 96938 254866 97174
rect 255102 96938 274546 97174
rect 274782 96938 274866 97174
rect 275102 96938 294546 97174
rect 294782 96938 294866 97174
rect 295102 96938 314546 97174
rect 314782 96938 314866 97174
rect 315102 96938 334546 97174
rect 334782 96938 334866 97174
rect 335102 96938 354546 97174
rect 354782 96938 354866 97174
rect 355102 96938 374546 97174
rect 374782 96938 374866 97174
rect 375102 96938 394546 97174
rect 394782 96938 394866 97174
rect 395102 96938 414546 97174
rect 414782 96938 414866 97174
rect 415102 96938 434546 97174
rect 434782 96938 434866 97174
rect 435102 96938 454546 97174
rect 454782 96938 454866 97174
rect 455102 96938 474546 97174
rect 474782 96938 474866 97174
rect 475102 96938 494546 97174
rect 494782 96938 494866 97174
rect 495102 96938 514546 97174
rect 514782 96938 514866 97174
rect 515102 96938 534546 97174
rect 534782 96938 534866 97174
rect 535102 96938 554546 97174
rect 554782 96938 554866 97174
rect 555102 96938 574546 97174
rect 574782 96938 574866 97174
rect 575102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 14546 96854
rect 14782 96618 14866 96854
rect 15102 96618 34546 96854
rect 34782 96618 34866 96854
rect 35102 96618 54546 96854
rect 54782 96618 54866 96854
rect 55102 96618 74546 96854
rect 74782 96618 74866 96854
rect 75102 96618 94546 96854
rect 94782 96618 94866 96854
rect 95102 96618 114546 96854
rect 114782 96618 114866 96854
rect 115102 96618 134546 96854
rect 134782 96618 134866 96854
rect 135102 96618 154546 96854
rect 154782 96618 154866 96854
rect 155102 96618 174546 96854
rect 174782 96618 174866 96854
rect 175102 96618 194546 96854
rect 194782 96618 194866 96854
rect 195102 96618 214546 96854
rect 214782 96618 214866 96854
rect 215102 96618 234546 96854
rect 234782 96618 234866 96854
rect 235102 96618 254546 96854
rect 254782 96618 254866 96854
rect 255102 96618 274546 96854
rect 274782 96618 274866 96854
rect 275102 96618 294546 96854
rect 294782 96618 294866 96854
rect 295102 96618 314546 96854
rect 314782 96618 314866 96854
rect 315102 96618 334546 96854
rect 334782 96618 334866 96854
rect 335102 96618 354546 96854
rect 354782 96618 354866 96854
rect 355102 96618 374546 96854
rect 374782 96618 374866 96854
rect 375102 96618 394546 96854
rect 394782 96618 394866 96854
rect 395102 96618 414546 96854
rect 414782 96618 414866 96854
rect 415102 96618 434546 96854
rect 434782 96618 434866 96854
rect 435102 96618 454546 96854
rect 454782 96618 454866 96854
rect 455102 96618 474546 96854
rect 474782 96618 474866 96854
rect 475102 96618 494546 96854
rect 494782 96618 494866 96854
rect 495102 96618 514546 96854
rect 514782 96618 514866 96854
rect 515102 96618 534546 96854
rect 534782 96618 534866 96854
rect 535102 96618 554546 96854
rect 554782 96618 554866 96854
rect 555102 96618 574546 96854
rect 574782 96618 574866 96854
rect 575102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 10826 93454
rect 11062 93218 11146 93454
rect 11382 93218 30826 93454
rect 31062 93218 31146 93454
rect 31382 93218 50826 93454
rect 51062 93218 51146 93454
rect 51382 93218 70826 93454
rect 71062 93218 71146 93454
rect 71382 93218 90826 93454
rect 91062 93218 91146 93454
rect 91382 93218 110826 93454
rect 111062 93218 111146 93454
rect 111382 93218 130826 93454
rect 131062 93218 131146 93454
rect 131382 93218 150826 93454
rect 151062 93218 151146 93454
rect 151382 93218 170826 93454
rect 171062 93218 171146 93454
rect 171382 93218 190826 93454
rect 191062 93218 191146 93454
rect 191382 93218 210826 93454
rect 211062 93218 211146 93454
rect 211382 93218 230826 93454
rect 231062 93218 231146 93454
rect 231382 93218 250826 93454
rect 251062 93218 251146 93454
rect 251382 93218 270826 93454
rect 271062 93218 271146 93454
rect 271382 93218 290826 93454
rect 291062 93218 291146 93454
rect 291382 93218 310826 93454
rect 311062 93218 311146 93454
rect 311382 93218 330826 93454
rect 331062 93218 331146 93454
rect 331382 93218 350826 93454
rect 351062 93218 351146 93454
rect 351382 93218 370826 93454
rect 371062 93218 371146 93454
rect 371382 93218 390826 93454
rect 391062 93218 391146 93454
rect 391382 93218 410826 93454
rect 411062 93218 411146 93454
rect 411382 93218 430826 93454
rect 431062 93218 431146 93454
rect 431382 93218 450826 93454
rect 451062 93218 451146 93454
rect 451382 93218 470826 93454
rect 471062 93218 471146 93454
rect 471382 93218 490826 93454
rect 491062 93218 491146 93454
rect 491382 93218 510826 93454
rect 511062 93218 511146 93454
rect 511382 93218 530826 93454
rect 531062 93218 531146 93454
rect 531382 93218 550826 93454
rect 551062 93218 551146 93454
rect 551382 93218 570826 93454
rect 571062 93218 571146 93454
rect 571382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 10826 93134
rect 11062 92898 11146 93134
rect 11382 92898 30826 93134
rect 31062 92898 31146 93134
rect 31382 92898 50826 93134
rect 51062 92898 51146 93134
rect 51382 92898 70826 93134
rect 71062 92898 71146 93134
rect 71382 92898 90826 93134
rect 91062 92898 91146 93134
rect 91382 92898 110826 93134
rect 111062 92898 111146 93134
rect 111382 92898 130826 93134
rect 131062 92898 131146 93134
rect 131382 92898 150826 93134
rect 151062 92898 151146 93134
rect 151382 92898 170826 93134
rect 171062 92898 171146 93134
rect 171382 92898 190826 93134
rect 191062 92898 191146 93134
rect 191382 92898 210826 93134
rect 211062 92898 211146 93134
rect 211382 92898 230826 93134
rect 231062 92898 231146 93134
rect 231382 92898 250826 93134
rect 251062 92898 251146 93134
rect 251382 92898 270826 93134
rect 271062 92898 271146 93134
rect 271382 92898 290826 93134
rect 291062 92898 291146 93134
rect 291382 92898 310826 93134
rect 311062 92898 311146 93134
rect 311382 92898 330826 93134
rect 331062 92898 331146 93134
rect 331382 92898 350826 93134
rect 351062 92898 351146 93134
rect 351382 92898 370826 93134
rect 371062 92898 371146 93134
rect 371382 92898 390826 93134
rect 391062 92898 391146 93134
rect 391382 92898 410826 93134
rect 411062 92898 411146 93134
rect 411382 92898 430826 93134
rect 431062 92898 431146 93134
rect 431382 92898 450826 93134
rect 451062 92898 451146 93134
rect 451382 92898 470826 93134
rect 471062 92898 471146 93134
rect 471382 92898 490826 93134
rect 491062 92898 491146 93134
rect 491382 92898 510826 93134
rect 511062 92898 511146 93134
rect 511382 92898 530826 93134
rect 531062 92898 531146 93134
rect 531382 92898 550826 93134
rect 551062 92898 551146 93134
rect 551382 92898 570826 93134
rect 571062 92898 571146 93134
rect 571382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 11986 86614
rect 12222 86378 12306 86614
rect 12542 86378 31986 86614
rect 32222 86378 32306 86614
rect 32542 86378 51986 86614
rect 52222 86378 52306 86614
rect 52542 86378 71986 86614
rect 72222 86378 72306 86614
rect 72542 86378 91986 86614
rect 92222 86378 92306 86614
rect 92542 86378 111986 86614
rect 112222 86378 112306 86614
rect 112542 86378 131986 86614
rect 132222 86378 132306 86614
rect 132542 86378 151986 86614
rect 152222 86378 152306 86614
rect 152542 86378 171986 86614
rect 172222 86378 172306 86614
rect 172542 86378 191986 86614
rect 192222 86378 192306 86614
rect 192542 86378 211986 86614
rect 212222 86378 212306 86614
rect 212542 86378 231986 86614
rect 232222 86378 232306 86614
rect 232542 86378 251986 86614
rect 252222 86378 252306 86614
rect 252542 86378 271986 86614
rect 272222 86378 272306 86614
rect 272542 86378 291986 86614
rect 292222 86378 292306 86614
rect 292542 86378 311986 86614
rect 312222 86378 312306 86614
rect 312542 86378 331986 86614
rect 332222 86378 332306 86614
rect 332542 86378 351986 86614
rect 352222 86378 352306 86614
rect 352542 86378 371986 86614
rect 372222 86378 372306 86614
rect 372542 86378 391986 86614
rect 392222 86378 392306 86614
rect 392542 86378 411986 86614
rect 412222 86378 412306 86614
rect 412542 86378 431986 86614
rect 432222 86378 432306 86614
rect 432542 86378 451986 86614
rect 452222 86378 452306 86614
rect 452542 86378 471986 86614
rect 472222 86378 472306 86614
rect 472542 86378 491986 86614
rect 492222 86378 492306 86614
rect 492542 86378 511986 86614
rect 512222 86378 512306 86614
rect 512542 86378 531986 86614
rect 532222 86378 532306 86614
rect 532542 86378 551986 86614
rect 552222 86378 552306 86614
rect 552542 86378 571986 86614
rect 572222 86378 572306 86614
rect 572542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 11986 86294
rect 12222 86058 12306 86294
rect 12542 86058 31986 86294
rect 32222 86058 32306 86294
rect 32542 86058 51986 86294
rect 52222 86058 52306 86294
rect 52542 86058 71986 86294
rect 72222 86058 72306 86294
rect 72542 86058 91986 86294
rect 92222 86058 92306 86294
rect 92542 86058 111986 86294
rect 112222 86058 112306 86294
rect 112542 86058 131986 86294
rect 132222 86058 132306 86294
rect 132542 86058 151986 86294
rect 152222 86058 152306 86294
rect 152542 86058 171986 86294
rect 172222 86058 172306 86294
rect 172542 86058 191986 86294
rect 192222 86058 192306 86294
rect 192542 86058 211986 86294
rect 212222 86058 212306 86294
rect 212542 86058 231986 86294
rect 232222 86058 232306 86294
rect 232542 86058 251986 86294
rect 252222 86058 252306 86294
rect 252542 86058 271986 86294
rect 272222 86058 272306 86294
rect 272542 86058 291986 86294
rect 292222 86058 292306 86294
rect 292542 86058 311986 86294
rect 312222 86058 312306 86294
rect 312542 86058 331986 86294
rect 332222 86058 332306 86294
rect 332542 86058 351986 86294
rect 352222 86058 352306 86294
rect 352542 86058 371986 86294
rect 372222 86058 372306 86294
rect 372542 86058 391986 86294
rect 392222 86058 392306 86294
rect 392542 86058 411986 86294
rect 412222 86058 412306 86294
rect 412542 86058 431986 86294
rect 432222 86058 432306 86294
rect 432542 86058 451986 86294
rect 452222 86058 452306 86294
rect 452542 86058 471986 86294
rect 472222 86058 472306 86294
rect 472542 86058 491986 86294
rect 492222 86058 492306 86294
rect 492542 86058 511986 86294
rect 512222 86058 512306 86294
rect 512542 86058 531986 86294
rect 532222 86058 532306 86294
rect 532542 86058 551986 86294
rect 552222 86058 552306 86294
rect 552542 86058 571986 86294
rect 572222 86058 572306 86294
rect 572542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 8266 82894
rect 8502 82658 8586 82894
rect 8822 82658 28266 82894
rect 28502 82658 28586 82894
rect 28822 82658 48266 82894
rect 48502 82658 48586 82894
rect 48822 82658 68266 82894
rect 68502 82658 68586 82894
rect 68822 82658 88266 82894
rect 88502 82658 88586 82894
rect 88822 82658 108266 82894
rect 108502 82658 108586 82894
rect 108822 82658 128266 82894
rect 128502 82658 128586 82894
rect 128822 82658 148266 82894
rect 148502 82658 148586 82894
rect 148822 82658 168266 82894
rect 168502 82658 168586 82894
rect 168822 82658 188266 82894
rect 188502 82658 188586 82894
rect 188822 82658 208266 82894
rect 208502 82658 208586 82894
rect 208822 82658 228266 82894
rect 228502 82658 228586 82894
rect 228822 82658 248266 82894
rect 248502 82658 248586 82894
rect 248822 82658 268266 82894
rect 268502 82658 268586 82894
rect 268822 82658 288266 82894
rect 288502 82658 288586 82894
rect 288822 82658 308266 82894
rect 308502 82658 308586 82894
rect 308822 82658 328266 82894
rect 328502 82658 328586 82894
rect 328822 82658 348266 82894
rect 348502 82658 348586 82894
rect 348822 82658 368266 82894
rect 368502 82658 368586 82894
rect 368822 82658 388266 82894
rect 388502 82658 388586 82894
rect 388822 82658 408266 82894
rect 408502 82658 408586 82894
rect 408822 82658 428266 82894
rect 428502 82658 428586 82894
rect 428822 82658 448266 82894
rect 448502 82658 448586 82894
rect 448822 82658 468266 82894
rect 468502 82658 468586 82894
rect 468822 82658 488266 82894
rect 488502 82658 488586 82894
rect 488822 82658 508266 82894
rect 508502 82658 508586 82894
rect 508822 82658 528266 82894
rect 528502 82658 528586 82894
rect 528822 82658 548266 82894
rect 548502 82658 548586 82894
rect 548822 82658 568266 82894
rect 568502 82658 568586 82894
rect 568822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 8266 82574
rect 8502 82338 8586 82574
rect 8822 82338 28266 82574
rect 28502 82338 28586 82574
rect 28822 82338 48266 82574
rect 48502 82338 48586 82574
rect 48822 82338 68266 82574
rect 68502 82338 68586 82574
rect 68822 82338 88266 82574
rect 88502 82338 88586 82574
rect 88822 82338 108266 82574
rect 108502 82338 108586 82574
rect 108822 82338 128266 82574
rect 128502 82338 128586 82574
rect 128822 82338 148266 82574
rect 148502 82338 148586 82574
rect 148822 82338 168266 82574
rect 168502 82338 168586 82574
rect 168822 82338 188266 82574
rect 188502 82338 188586 82574
rect 188822 82338 208266 82574
rect 208502 82338 208586 82574
rect 208822 82338 228266 82574
rect 228502 82338 228586 82574
rect 228822 82338 248266 82574
rect 248502 82338 248586 82574
rect 248822 82338 268266 82574
rect 268502 82338 268586 82574
rect 268822 82338 288266 82574
rect 288502 82338 288586 82574
rect 288822 82338 308266 82574
rect 308502 82338 308586 82574
rect 308822 82338 328266 82574
rect 328502 82338 328586 82574
rect 328822 82338 348266 82574
rect 348502 82338 348586 82574
rect 348822 82338 368266 82574
rect 368502 82338 368586 82574
rect 368822 82338 388266 82574
rect 388502 82338 388586 82574
rect 388822 82338 408266 82574
rect 408502 82338 408586 82574
rect 408822 82338 428266 82574
rect 428502 82338 428586 82574
rect 428822 82338 448266 82574
rect 448502 82338 448586 82574
rect 448822 82338 468266 82574
rect 468502 82338 468586 82574
rect 468822 82338 488266 82574
rect 488502 82338 488586 82574
rect 488822 82338 508266 82574
rect 508502 82338 508586 82574
rect 508822 82338 528266 82574
rect 528502 82338 528586 82574
rect 528822 82338 548266 82574
rect 548502 82338 548586 82574
rect 548822 82338 568266 82574
rect 568502 82338 568586 82574
rect 568822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 4546 79174
rect 4782 78938 4866 79174
rect 5102 78938 24546 79174
rect 24782 78938 24866 79174
rect 25102 78938 44546 79174
rect 44782 78938 44866 79174
rect 45102 78938 64546 79174
rect 64782 78938 64866 79174
rect 65102 78938 84546 79174
rect 84782 78938 84866 79174
rect 85102 78938 104546 79174
rect 104782 78938 104866 79174
rect 105102 78938 124546 79174
rect 124782 78938 124866 79174
rect 125102 78938 144546 79174
rect 144782 78938 144866 79174
rect 145102 78938 164546 79174
rect 164782 78938 164866 79174
rect 165102 78938 184546 79174
rect 184782 78938 184866 79174
rect 185102 78938 204546 79174
rect 204782 78938 204866 79174
rect 205102 78938 224546 79174
rect 224782 78938 224866 79174
rect 225102 78938 244546 79174
rect 244782 78938 244866 79174
rect 245102 78938 264546 79174
rect 264782 78938 264866 79174
rect 265102 78938 284546 79174
rect 284782 78938 284866 79174
rect 285102 78938 304546 79174
rect 304782 78938 304866 79174
rect 305102 78938 324546 79174
rect 324782 78938 324866 79174
rect 325102 78938 344546 79174
rect 344782 78938 344866 79174
rect 345102 78938 364546 79174
rect 364782 78938 364866 79174
rect 365102 78938 384546 79174
rect 384782 78938 384866 79174
rect 385102 78938 404546 79174
rect 404782 78938 404866 79174
rect 405102 78938 424546 79174
rect 424782 78938 424866 79174
rect 425102 78938 444546 79174
rect 444782 78938 444866 79174
rect 445102 78938 464546 79174
rect 464782 78938 464866 79174
rect 465102 78938 484546 79174
rect 484782 78938 484866 79174
rect 485102 78938 504546 79174
rect 504782 78938 504866 79174
rect 505102 78938 524546 79174
rect 524782 78938 524866 79174
rect 525102 78938 544546 79174
rect 544782 78938 544866 79174
rect 545102 78938 564546 79174
rect 564782 78938 564866 79174
rect 565102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 4546 78854
rect 4782 78618 4866 78854
rect 5102 78618 24546 78854
rect 24782 78618 24866 78854
rect 25102 78618 44546 78854
rect 44782 78618 44866 78854
rect 45102 78618 64546 78854
rect 64782 78618 64866 78854
rect 65102 78618 84546 78854
rect 84782 78618 84866 78854
rect 85102 78618 104546 78854
rect 104782 78618 104866 78854
rect 105102 78618 124546 78854
rect 124782 78618 124866 78854
rect 125102 78618 144546 78854
rect 144782 78618 144866 78854
rect 145102 78618 164546 78854
rect 164782 78618 164866 78854
rect 165102 78618 184546 78854
rect 184782 78618 184866 78854
rect 185102 78618 204546 78854
rect 204782 78618 204866 78854
rect 205102 78618 224546 78854
rect 224782 78618 224866 78854
rect 225102 78618 244546 78854
rect 244782 78618 244866 78854
rect 245102 78618 264546 78854
rect 264782 78618 264866 78854
rect 265102 78618 284546 78854
rect 284782 78618 284866 78854
rect 285102 78618 304546 78854
rect 304782 78618 304866 78854
rect 305102 78618 324546 78854
rect 324782 78618 324866 78854
rect 325102 78618 344546 78854
rect 344782 78618 344866 78854
rect 345102 78618 364546 78854
rect 364782 78618 364866 78854
rect 365102 78618 384546 78854
rect 384782 78618 384866 78854
rect 385102 78618 404546 78854
rect 404782 78618 404866 78854
rect 405102 78618 424546 78854
rect 424782 78618 424866 78854
rect 425102 78618 444546 78854
rect 444782 78618 444866 78854
rect 445102 78618 464546 78854
rect 464782 78618 464866 78854
rect 465102 78618 484546 78854
rect 484782 78618 484866 78854
rect 485102 78618 504546 78854
rect 504782 78618 504866 78854
rect 505102 78618 524546 78854
rect 524782 78618 524866 78854
rect 525102 78618 544546 78854
rect 544782 78618 544866 78854
rect 545102 78618 564546 78854
rect 564782 78618 564866 78854
rect 565102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 826 75454
rect 1062 75218 1146 75454
rect 1382 75218 20826 75454
rect 21062 75218 21146 75454
rect 21382 75218 40826 75454
rect 41062 75218 41146 75454
rect 41382 75218 60826 75454
rect 61062 75218 61146 75454
rect 61382 75218 80826 75454
rect 81062 75218 81146 75454
rect 81382 75218 100826 75454
rect 101062 75218 101146 75454
rect 101382 75218 120826 75454
rect 121062 75218 121146 75454
rect 121382 75218 140826 75454
rect 141062 75218 141146 75454
rect 141382 75218 160826 75454
rect 161062 75218 161146 75454
rect 161382 75218 180826 75454
rect 181062 75218 181146 75454
rect 181382 75218 200826 75454
rect 201062 75218 201146 75454
rect 201382 75218 220826 75454
rect 221062 75218 221146 75454
rect 221382 75218 240826 75454
rect 241062 75218 241146 75454
rect 241382 75218 260826 75454
rect 261062 75218 261146 75454
rect 261382 75218 280826 75454
rect 281062 75218 281146 75454
rect 281382 75218 300826 75454
rect 301062 75218 301146 75454
rect 301382 75218 320826 75454
rect 321062 75218 321146 75454
rect 321382 75218 340826 75454
rect 341062 75218 341146 75454
rect 341382 75218 360826 75454
rect 361062 75218 361146 75454
rect 361382 75218 380826 75454
rect 381062 75218 381146 75454
rect 381382 75218 400826 75454
rect 401062 75218 401146 75454
rect 401382 75218 420826 75454
rect 421062 75218 421146 75454
rect 421382 75218 440826 75454
rect 441062 75218 441146 75454
rect 441382 75218 460826 75454
rect 461062 75218 461146 75454
rect 461382 75218 480826 75454
rect 481062 75218 481146 75454
rect 481382 75218 500826 75454
rect 501062 75218 501146 75454
rect 501382 75218 520826 75454
rect 521062 75218 521146 75454
rect 521382 75218 540826 75454
rect 541062 75218 541146 75454
rect 541382 75218 560826 75454
rect 561062 75218 561146 75454
rect 561382 75218 580826 75454
rect 581062 75218 581146 75454
rect 581382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 826 75134
rect 1062 74898 1146 75134
rect 1382 74898 20826 75134
rect 21062 74898 21146 75134
rect 21382 74898 40826 75134
rect 41062 74898 41146 75134
rect 41382 74898 60826 75134
rect 61062 74898 61146 75134
rect 61382 74898 80826 75134
rect 81062 74898 81146 75134
rect 81382 74898 100826 75134
rect 101062 74898 101146 75134
rect 101382 74898 120826 75134
rect 121062 74898 121146 75134
rect 121382 74898 140826 75134
rect 141062 74898 141146 75134
rect 141382 74898 160826 75134
rect 161062 74898 161146 75134
rect 161382 74898 180826 75134
rect 181062 74898 181146 75134
rect 181382 74898 200826 75134
rect 201062 74898 201146 75134
rect 201382 74898 220826 75134
rect 221062 74898 221146 75134
rect 221382 74898 240826 75134
rect 241062 74898 241146 75134
rect 241382 74898 260826 75134
rect 261062 74898 261146 75134
rect 261382 74898 280826 75134
rect 281062 74898 281146 75134
rect 281382 74898 300826 75134
rect 301062 74898 301146 75134
rect 301382 74898 320826 75134
rect 321062 74898 321146 75134
rect 321382 74898 340826 75134
rect 341062 74898 341146 75134
rect 341382 74898 360826 75134
rect 361062 74898 361146 75134
rect 361382 74898 380826 75134
rect 381062 74898 381146 75134
rect 381382 74898 400826 75134
rect 401062 74898 401146 75134
rect 401382 74898 420826 75134
rect 421062 74898 421146 75134
rect 421382 74898 440826 75134
rect 441062 74898 441146 75134
rect 441382 74898 460826 75134
rect 461062 74898 461146 75134
rect 461382 74898 480826 75134
rect 481062 74898 481146 75134
rect 481382 74898 500826 75134
rect 501062 74898 501146 75134
rect 501382 74898 520826 75134
rect 521062 74898 521146 75134
rect 521382 74898 540826 75134
rect 541062 74898 541146 75134
rect 541382 74898 560826 75134
rect 561062 74898 561146 75134
rect 561382 74898 580826 75134
rect 581062 74898 581146 75134
rect 581382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 81986 68614
rect 82222 68378 82306 68614
rect 82542 68378 101986 68614
rect 102222 68378 102306 68614
rect 102542 68378 121986 68614
rect 122222 68378 122306 68614
rect 122542 68378 141986 68614
rect 142222 68378 142306 68614
rect 142542 68378 161986 68614
rect 162222 68378 162306 68614
rect 162542 68378 181986 68614
rect 182222 68378 182306 68614
rect 182542 68378 201986 68614
rect 202222 68378 202306 68614
rect 202542 68378 221986 68614
rect 222222 68378 222306 68614
rect 222542 68378 241986 68614
rect 242222 68378 242306 68614
rect 242542 68378 261986 68614
rect 262222 68378 262306 68614
rect 262542 68378 281986 68614
rect 282222 68378 282306 68614
rect 282542 68378 301986 68614
rect 302222 68378 302306 68614
rect 302542 68378 321986 68614
rect 322222 68378 322306 68614
rect 322542 68378 341986 68614
rect 342222 68378 342306 68614
rect 342542 68378 361986 68614
rect 362222 68378 362306 68614
rect 362542 68378 381986 68614
rect 382222 68378 382306 68614
rect 382542 68378 401986 68614
rect 402222 68378 402306 68614
rect 402542 68378 421986 68614
rect 422222 68378 422306 68614
rect 422542 68378 441986 68614
rect 442222 68378 442306 68614
rect 442542 68378 461986 68614
rect 462222 68378 462306 68614
rect 462542 68378 481986 68614
rect 482222 68378 482306 68614
rect 482542 68378 501986 68614
rect 502222 68378 502306 68614
rect 502542 68378 521986 68614
rect 522222 68378 522306 68614
rect 522542 68378 541986 68614
rect 542222 68378 542306 68614
rect 542542 68378 561986 68614
rect 562222 68378 562306 68614
rect 562542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 81986 68294
rect 82222 68058 82306 68294
rect 82542 68058 101986 68294
rect 102222 68058 102306 68294
rect 102542 68058 121986 68294
rect 122222 68058 122306 68294
rect 122542 68058 141986 68294
rect 142222 68058 142306 68294
rect 142542 68058 161986 68294
rect 162222 68058 162306 68294
rect 162542 68058 181986 68294
rect 182222 68058 182306 68294
rect 182542 68058 201986 68294
rect 202222 68058 202306 68294
rect 202542 68058 221986 68294
rect 222222 68058 222306 68294
rect 222542 68058 241986 68294
rect 242222 68058 242306 68294
rect 242542 68058 261986 68294
rect 262222 68058 262306 68294
rect 262542 68058 281986 68294
rect 282222 68058 282306 68294
rect 282542 68058 301986 68294
rect 302222 68058 302306 68294
rect 302542 68058 321986 68294
rect 322222 68058 322306 68294
rect 322542 68058 341986 68294
rect 342222 68058 342306 68294
rect 342542 68058 361986 68294
rect 362222 68058 362306 68294
rect 362542 68058 381986 68294
rect 382222 68058 382306 68294
rect 382542 68058 401986 68294
rect 402222 68058 402306 68294
rect 402542 68058 421986 68294
rect 422222 68058 422306 68294
rect 422542 68058 441986 68294
rect 442222 68058 442306 68294
rect 442542 68058 461986 68294
rect 462222 68058 462306 68294
rect 462542 68058 481986 68294
rect 482222 68058 482306 68294
rect 482542 68058 501986 68294
rect 502222 68058 502306 68294
rect 502542 68058 521986 68294
rect 522222 68058 522306 68294
rect 522542 68058 541986 68294
rect 542222 68058 542306 68294
rect 542542 68058 561986 68294
rect 562222 68058 562306 68294
rect 562542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 78266 64894
rect 78502 64658 78586 64894
rect 78822 64658 98266 64894
rect 98502 64658 98586 64894
rect 98822 64658 118266 64894
rect 118502 64658 118586 64894
rect 118822 64658 138266 64894
rect 138502 64658 138586 64894
rect 138822 64658 158266 64894
rect 158502 64658 158586 64894
rect 158822 64658 178266 64894
rect 178502 64658 178586 64894
rect 178822 64658 198266 64894
rect 198502 64658 198586 64894
rect 198822 64658 218266 64894
rect 218502 64658 218586 64894
rect 218822 64658 238266 64894
rect 238502 64658 238586 64894
rect 238822 64658 258266 64894
rect 258502 64658 258586 64894
rect 258822 64658 278266 64894
rect 278502 64658 278586 64894
rect 278822 64658 298266 64894
rect 298502 64658 298586 64894
rect 298822 64658 318266 64894
rect 318502 64658 318586 64894
rect 318822 64658 338266 64894
rect 338502 64658 338586 64894
rect 338822 64658 358266 64894
rect 358502 64658 358586 64894
rect 358822 64658 378266 64894
rect 378502 64658 378586 64894
rect 378822 64658 398266 64894
rect 398502 64658 398586 64894
rect 398822 64658 418266 64894
rect 418502 64658 418586 64894
rect 418822 64658 438266 64894
rect 438502 64658 438586 64894
rect 438822 64658 458266 64894
rect 458502 64658 458586 64894
rect 458822 64658 478266 64894
rect 478502 64658 478586 64894
rect 478822 64658 498266 64894
rect 498502 64658 498586 64894
rect 498822 64658 518266 64894
rect 518502 64658 518586 64894
rect 518822 64658 538266 64894
rect 538502 64658 538586 64894
rect 538822 64658 558266 64894
rect 558502 64658 558586 64894
rect 558822 64658 578266 64894
rect 578502 64658 578586 64894
rect 578822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 78266 64574
rect 78502 64338 78586 64574
rect 78822 64338 98266 64574
rect 98502 64338 98586 64574
rect 98822 64338 118266 64574
rect 118502 64338 118586 64574
rect 118822 64338 138266 64574
rect 138502 64338 138586 64574
rect 138822 64338 158266 64574
rect 158502 64338 158586 64574
rect 158822 64338 178266 64574
rect 178502 64338 178586 64574
rect 178822 64338 198266 64574
rect 198502 64338 198586 64574
rect 198822 64338 218266 64574
rect 218502 64338 218586 64574
rect 218822 64338 238266 64574
rect 238502 64338 238586 64574
rect 238822 64338 258266 64574
rect 258502 64338 258586 64574
rect 258822 64338 278266 64574
rect 278502 64338 278586 64574
rect 278822 64338 298266 64574
rect 298502 64338 298586 64574
rect 298822 64338 318266 64574
rect 318502 64338 318586 64574
rect 318822 64338 338266 64574
rect 338502 64338 338586 64574
rect 338822 64338 358266 64574
rect 358502 64338 358586 64574
rect 358822 64338 378266 64574
rect 378502 64338 378586 64574
rect 378822 64338 398266 64574
rect 398502 64338 398586 64574
rect 398822 64338 418266 64574
rect 418502 64338 418586 64574
rect 418822 64338 438266 64574
rect 438502 64338 438586 64574
rect 438822 64338 458266 64574
rect 458502 64338 458586 64574
rect 458822 64338 478266 64574
rect 478502 64338 478586 64574
rect 478822 64338 498266 64574
rect 498502 64338 498586 64574
rect 498822 64338 518266 64574
rect 518502 64338 518586 64574
rect 518822 64338 538266 64574
rect 538502 64338 538586 64574
rect 538822 64338 558266 64574
rect 558502 64338 558586 64574
rect 558822 64338 578266 64574
rect 578502 64338 578586 64574
rect 578822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 14546 61174
rect 14782 60938 14866 61174
rect 15102 60938 74546 61174
rect 74782 60938 74866 61174
rect 75102 60938 94546 61174
rect 94782 60938 94866 61174
rect 95102 60938 114546 61174
rect 114782 60938 114866 61174
rect 115102 60938 134546 61174
rect 134782 60938 134866 61174
rect 135102 60938 154546 61174
rect 154782 60938 154866 61174
rect 155102 60938 174546 61174
rect 174782 60938 174866 61174
rect 175102 60938 194546 61174
rect 194782 60938 194866 61174
rect 195102 60938 214546 61174
rect 214782 60938 214866 61174
rect 215102 60938 234546 61174
rect 234782 60938 234866 61174
rect 235102 60938 254546 61174
rect 254782 60938 254866 61174
rect 255102 60938 274546 61174
rect 274782 60938 274866 61174
rect 275102 60938 294546 61174
rect 294782 60938 294866 61174
rect 295102 60938 314546 61174
rect 314782 60938 314866 61174
rect 315102 60938 334546 61174
rect 334782 60938 334866 61174
rect 335102 60938 354546 61174
rect 354782 60938 354866 61174
rect 355102 60938 374546 61174
rect 374782 60938 374866 61174
rect 375102 60938 394546 61174
rect 394782 60938 394866 61174
rect 395102 60938 414546 61174
rect 414782 60938 414866 61174
rect 415102 60938 434546 61174
rect 434782 60938 434866 61174
rect 435102 60938 454546 61174
rect 454782 60938 454866 61174
rect 455102 60938 474546 61174
rect 474782 60938 474866 61174
rect 475102 60938 494546 61174
rect 494782 60938 494866 61174
rect 495102 60938 514546 61174
rect 514782 60938 514866 61174
rect 515102 60938 534546 61174
rect 534782 60938 534866 61174
rect 535102 60938 554546 61174
rect 554782 60938 554866 61174
rect 555102 60938 574546 61174
rect 574782 60938 574866 61174
rect 575102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 14546 60854
rect 14782 60618 14866 60854
rect 15102 60618 74546 60854
rect 74782 60618 74866 60854
rect 75102 60618 94546 60854
rect 94782 60618 94866 60854
rect 95102 60618 114546 60854
rect 114782 60618 114866 60854
rect 115102 60618 134546 60854
rect 134782 60618 134866 60854
rect 135102 60618 154546 60854
rect 154782 60618 154866 60854
rect 155102 60618 174546 60854
rect 174782 60618 174866 60854
rect 175102 60618 194546 60854
rect 194782 60618 194866 60854
rect 195102 60618 214546 60854
rect 214782 60618 214866 60854
rect 215102 60618 234546 60854
rect 234782 60618 234866 60854
rect 235102 60618 254546 60854
rect 254782 60618 254866 60854
rect 255102 60618 274546 60854
rect 274782 60618 274866 60854
rect 275102 60618 294546 60854
rect 294782 60618 294866 60854
rect 295102 60618 314546 60854
rect 314782 60618 314866 60854
rect 315102 60618 334546 60854
rect 334782 60618 334866 60854
rect 335102 60618 354546 60854
rect 354782 60618 354866 60854
rect 355102 60618 374546 60854
rect 374782 60618 374866 60854
rect 375102 60618 394546 60854
rect 394782 60618 394866 60854
rect 395102 60618 414546 60854
rect 414782 60618 414866 60854
rect 415102 60618 434546 60854
rect 434782 60618 434866 60854
rect 435102 60618 454546 60854
rect 454782 60618 454866 60854
rect 455102 60618 474546 60854
rect 474782 60618 474866 60854
rect 475102 60618 494546 60854
rect 494782 60618 494866 60854
rect 495102 60618 514546 60854
rect 514782 60618 514866 60854
rect 515102 60618 534546 60854
rect 534782 60618 534866 60854
rect 535102 60618 554546 60854
rect 554782 60618 554866 60854
rect 555102 60618 574546 60854
rect 574782 60618 574866 60854
rect 575102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 10826 57454
rect 11062 57218 11146 57454
rect 11382 57218 39610 57454
rect 39846 57218 90826 57454
rect 91062 57218 91146 57454
rect 91382 57218 110826 57454
rect 111062 57218 111146 57454
rect 111382 57218 130826 57454
rect 131062 57218 131146 57454
rect 131382 57218 150826 57454
rect 151062 57218 151146 57454
rect 151382 57218 170826 57454
rect 171062 57218 171146 57454
rect 171382 57218 190826 57454
rect 191062 57218 191146 57454
rect 191382 57218 210826 57454
rect 211062 57218 211146 57454
rect 211382 57218 230826 57454
rect 231062 57218 231146 57454
rect 231382 57218 250826 57454
rect 251062 57218 251146 57454
rect 251382 57218 270826 57454
rect 271062 57218 271146 57454
rect 271382 57218 290826 57454
rect 291062 57218 291146 57454
rect 291382 57218 310826 57454
rect 311062 57218 311146 57454
rect 311382 57218 330826 57454
rect 331062 57218 331146 57454
rect 331382 57218 350826 57454
rect 351062 57218 351146 57454
rect 351382 57218 370826 57454
rect 371062 57218 371146 57454
rect 371382 57218 390826 57454
rect 391062 57218 391146 57454
rect 391382 57218 410826 57454
rect 411062 57218 411146 57454
rect 411382 57218 430826 57454
rect 431062 57218 431146 57454
rect 431382 57218 450826 57454
rect 451062 57218 451146 57454
rect 451382 57218 470826 57454
rect 471062 57218 471146 57454
rect 471382 57218 490826 57454
rect 491062 57218 491146 57454
rect 491382 57218 510826 57454
rect 511062 57218 511146 57454
rect 511382 57218 530826 57454
rect 531062 57218 531146 57454
rect 531382 57218 550826 57454
rect 551062 57218 551146 57454
rect 551382 57218 570826 57454
rect 571062 57218 571146 57454
rect 571382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 10826 57134
rect 11062 56898 11146 57134
rect 11382 56898 39610 57134
rect 39846 56898 90826 57134
rect 91062 56898 91146 57134
rect 91382 56898 110826 57134
rect 111062 56898 111146 57134
rect 111382 56898 130826 57134
rect 131062 56898 131146 57134
rect 131382 56898 150826 57134
rect 151062 56898 151146 57134
rect 151382 56898 170826 57134
rect 171062 56898 171146 57134
rect 171382 56898 190826 57134
rect 191062 56898 191146 57134
rect 191382 56898 210826 57134
rect 211062 56898 211146 57134
rect 211382 56898 230826 57134
rect 231062 56898 231146 57134
rect 231382 56898 250826 57134
rect 251062 56898 251146 57134
rect 251382 56898 270826 57134
rect 271062 56898 271146 57134
rect 271382 56898 290826 57134
rect 291062 56898 291146 57134
rect 291382 56898 310826 57134
rect 311062 56898 311146 57134
rect 311382 56898 330826 57134
rect 331062 56898 331146 57134
rect 331382 56898 350826 57134
rect 351062 56898 351146 57134
rect 351382 56898 370826 57134
rect 371062 56898 371146 57134
rect 371382 56898 390826 57134
rect 391062 56898 391146 57134
rect 391382 56898 410826 57134
rect 411062 56898 411146 57134
rect 411382 56898 430826 57134
rect 431062 56898 431146 57134
rect 431382 56898 450826 57134
rect 451062 56898 451146 57134
rect 451382 56898 470826 57134
rect 471062 56898 471146 57134
rect 471382 56898 490826 57134
rect 491062 56898 491146 57134
rect 491382 56898 510826 57134
rect 511062 56898 511146 57134
rect 511382 56898 530826 57134
rect 531062 56898 531146 57134
rect 531382 56898 550826 57134
rect 551062 56898 551146 57134
rect 551382 56898 570826 57134
rect 571062 56898 571146 57134
rect 571382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 11986 50614
rect 12222 50378 12306 50614
rect 12542 50378 91986 50614
rect 92222 50378 92306 50614
rect 92542 50378 111986 50614
rect 112222 50378 112306 50614
rect 112542 50378 131986 50614
rect 132222 50378 132306 50614
rect 132542 50378 151986 50614
rect 152222 50378 152306 50614
rect 152542 50378 171986 50614
rect 172222 50378 172306 50614
rect 172542 50378 191986 50614
rect 192222 50378 192306 50614
rect 192542 50378 211986 50614
rect 212222 50378 212306 50614
rect 212542 50378 231986 50614
rect 232222 50378 232306 50614
rect 232542 50378 251986 50614
rect 252222 50378 252306 50614
rect 252542 50378 271986 50614
rect 272222 50378 272306 50614
rect 272542 50378 291986 50614
rect 292222 50378 292306 50614
rect 292542 50378 311986 50614
rect 312222 50378 312306 50614
rect 312542 50378 331986 50614
rect 332222 50378 332306 50614
rect 332542 50378 351986 50614
rect 352222 50378 352306 50614
rect 352542 50378 371986 50614
rect 372222 50378 372306 50614
rect 372542 50378 391986 50614
rect 392222 50378 392306 50614
rect 392542 50378 411986 50614
rect 412222 50378 412306 50614
rect 412542 50378 431986 50614
rect 432222 50378 432306 50614
rect 432542 50378 451986 50614
rect 452222 50378 452306 50614
rect 452542 50378 471986 50614
rect 472222 50378 472306 50614
rect 472542 50378 491986 50614
rect 492222 50378 492306 50614
rect 492542 50378 511986 50614
rect 512222 50378 512306 50614
rect 512542 50378 531986 50614
rect 532222 50378 532306 50614
rect 532542 50378 551986 50614
rect 552222 50378 552306 50614
rect 552542 50378 571986 50614
rect 572222 50378 572306 50614
rect 572542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 11986 50294
rect 12222 50058 12306 50294
rect 12542 50058 91986 50294
rect 92222 50058 92306 50294
rect 92542 50058 111986 50294
rect 112222 50058 112306 50294
rect 112542 50058 131986 50294
rect 132222 50058 132306 50294
rect 132542 50058 151986 50294
rect 152222 50058 152306 50294
rect 152542 50058 171986 50294
rect 172222 50058 172306 50294
rect 172542 50058 191986 50294
rect 192222 50058 192306 50294
rect 192542 50058 211986 50294
rect 212222 50058 212306 50294
rect 212542 50058 231986 50294
rect 232222 50058 232306 50294
rect 232542 50058 251986 50294
rect 252222 50058 252306 50294
rect 252542 50058 271986 50294
rect 272222 50058 272306 50294
rect 272542 50058 291986 50294
rect 292222 50058 292306 50294
rect 292542 50058 311986 50294
rect 312222 50058 312306 50294
rect 312542 50058 331986 50294
rect 332222 50058 332306 50294
rect 332542 50058 351986 50294
rect 352222 50058 352306 50294
rect 352542 50058 371986 50294
rect 372222 50058 372306 50294
rect 372542 50058 391986 50294
rect 392222 50058 392306 50294
rect 392542 50058 411986 50294
rect 412222 50058 412306 50294
rect 412542 50058 431986 50294
rect 432222 50058 432306 50294
rect 432542 50058 451986 50294
rect 452222 50058 452306 50294
rect 452542 50058 471986 50294
rect 472222 50058 472306 50294
rect 472542 50058 491986 50294
rect 492222 50058 492306 50294
rect 492542 50058 511986 50294
rect 512222 50058 512306 50294
rect 512542 50058 531986 50294
rect 532222 50058 532306 50294
rect 532542 50058 551986 50294
rect 552222 50058 552306 50294
rect 552542 50058 571986 50294
rect 572222 50058 572306 50294
rect 572542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 8266 46894
rect 8502 46658 8586 46894
rect 8822 46658 88266 46894
rect 88502 46658 88586 46894
rect 88822 46658 108266 46894
rect 108502 46658 108586 46894
rect 108822 46658 128266 46894
rect 128502 46658 128586 46894
rect 128822 46658 148266 46894
rect 148502 46658 148586 46894
rect 148822 46658 168266 46894
rect 168502 46658 168586 46894
rect 168822 46658 188266 46894
rect 188502 46658 188586 46894
rect 188822 46658 208266 46894
rect 208502 46658 208586 46894
rect 208822 46658 228266 46894
rect 228502 46658 228586 46894
rect 228822 46658 248266 46894
rect 248502 46658 248586 46894
rect 248822 46658 268266 46894
rect 268502 46658 268586 46894
rect 268822 46658 288266 46894
rect 288502 46658 288586 46894
rect 288822 46658 308266 46894
rect 308502 46658 308586 46894
rect 308822 46658 328266 46894
rect 328502 46658 328586 46894
rect 328822 46658 348266 46894
rect 348502 46658 348586 46894
rect 348822 46658 368266 46894
rect 368502 46658 368586 46894
rect 368822 46658 388266 46894
rect 388502 46658 388586 46894
rect 388822 46658 408266 46894
rect 408502 46658 408586 46894
rect 408822 46658 428266 46894
rect 428502 46658 428586 46894
rect 428822 46658 448266 46894
rect 448502 46658 448586 46894
rect 448822 46658 468266 46894
rect 468502 46658 468586 46894
rect 468822 46658 488266 46894
rect 488502 46658 488586 46894
rect 488822 46658 508266 46894
rect 508502 46658 508586 46894
rect 508822 46658 528266 46894
rect 528502 46658 528586 46894
rect 528822 46658 548266 46894
rect 548502 46658 548586 46894
rect 548822 46658 568266 46894
rect 568502 46658 568586 46894
rect 568822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 8266 46574
rect 8502 46338 8586 46574
rect 8822 46338 88266 46574
rect 88502 46338 88586 46574
rect 88822 46338 108266 46574
rect 108502 46338 108586 46574
rect 108822 46338 128266 46574
rect 128502 46338 128586 46574
rect 128822 46338 148266 46574
rect 148502 46338 148586 46574
rect 148822 46338 168266 46574
rect 168502 46338 168586 46574
rect 168822 46338 188266 46574
rect 188502 46338 188586 46574
rect 188822 46338 208266 46574
rect 208502 46338 208586 46574
rect 208822 46338 228266 46574
rect 228502 46338 228586 46574
rect 228822 46338 248266 46574
rect 248502 46338 248586 46574
rect 248822 46338 268266 46574
rect 268502 46338 268586 46574
rect 268822 46338 288266 46574
rect 288502 46338 288586 46574
rect 288822 46338 308266 46574
rect 308502 46338 308586 46574
rect 308822 46338 328266 46574
rect 328502 46338 328586 46574
rect 328822 46338 348266 46574
rect 348502 46338 348586 46574
rect 348822 46338 368266 46574
rect 368502 46338 368586 46574
rect 368822 46338 388266 46574
rect 388502 46338 388586 46574
rect 388822 46338 408266 46574
rect 408502 46338 408586 46574
rect 408822 46338 428266 46574
rect 428502 46338 428586 46574
rect 428822 46338 448266 46574
rect 448502 46338 448586 46574
rect 448822 46338 468266 46574
rect 468502 46338 468586 46574
rect 468822 46338 488266 46574
rect 488502 46338 488586 46574
rect 488822 46338 508266 46574
rect 508502 46338 508586 46574
rect 508822 46338 528266 46574
rect 528502 46338 528586 46574
rect 528822 46338 548266 46574
rect 548502 46338 548586 46574
rect 548822 46338 568266 46574
rect 568502 46338 568586 46574
rect 568822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 4546 43174
rect 4782 42938 4866 43174
rect 5102 42938 84546 43174
rect 84782 42938 84866 43174
rect 85102 42938 104546 43174
rect 104782 42938 104866 43174
rect 105102 42938 124546 43174
rect 124782 42938 124866 43174
rect 125102 42938 144546 43174
rect 144782 42938 144866 43174
rect 145102 42938 164546 43174
rect 164782 42938 164866 43174
rect 165102 42938 184546 43174
rect 184782 42938 184866 43174
rect 185102 42938 204546 43174
rect 204782 42938 204866 43174
rect 205102 42938 224546 43174
rect 224782 42938 224866 43174
rect 225102 42938 244546 43174
rect 244782 42938 244866 43174
rect 245102 42938 264546 43174
rect 264782 42938 264866 43174
rect 265102 42938 284546 43174
rect 284782 42938 284866 43174
rect 285102 42938 304546 43174
rect 304782 42938 304866 43174
rect 305102 42938 324546 43174
rect 324782 42938 324866 43174
rect 325102 42938 344546 43174
rect 344782 42938 344866 43174
rect 345102 42938 364546 43174
rect 364782 42938 364866 43174
rect 365102 42938 384546 43174
rect 384782 42938 384866 43174
rect 385102 42938 404546 43174
rect 404782 42938 404866 43174
rect 405102 42938 424546 43174
rect 424782 42938 424866 43174
rect 425102 42938 444546 43174
rect 444782 42938 444866 43174
rect 445102 42938 464546 43174
rect 464782 42938 464866 43174
rect 465102 42938 484546 43174
rect 484782 42938 484866 43174
rect 485102 42938 504546 43174
rect 504782 42938 504866 43174
rect 505102 42938 524546 43174
rect 524782 42938 524866 43174
rect 525102 42938 544546 43174
rect 544782 42938 544866 43174
rect 545102 42938 564546 43174
rect 564782 42938 564866 43174
rect 565102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 4546 42854
rect 4782 42618 4866 42854
rect 5102 42618 84546 42854
rect 84782 42618 84866 42854
rect 85102 42618 104546 42854
rect 104782 42618 104866 42854
rect 105102 42618 124546 42854
rect 124782 42618 124866 42854
rect 125102 42618 144546 42854
rect 144782 42618 144866 42854
rect 145102 42618 164546 42854
rect 164782 42618 164866 42854
rect 165102 42618 184546 42854
rect 184782 42618 184866 42854
rect 185102 42618 204546 42854
rect 204782 42618 204866 42854
rect 205102 42618 224546 42854
rect 224782 42618 224866 42854
rect 225102 42618 244546 42854
rect 244782 42618 244866 42854
rect 245102 42618 264546 42854
rect 264782 42618 264866 42854
rect 265102 42618 284546 42854
rect 284782 42618 284866 42854
rect 285102 42618 304546 42854
rect 304782 42618 304866 42854
rect 305102 42618 324546 42854
rect 324782 42618 324866 42854
rect 325102 42618 344546 42854
rect 344782 42618 344866 42854
rect 345102 42618 364546 42854
rect 364782 42618 364866 42854
rect 365102 42618 384546 42854
rect 384782 42618 384866 42854
rect 385102 42618 404546 42854
rect 404782 42618 404866 42854
rect 405102 42618 424546 42854
rect 424782 42618 424866 42854
rect 425102 42618 444546 42854
rect 444782 42618 444866 42854
rect 445102 42618 464546 42854
rect 464782 42618 464866 42854
rect 465102 42618 484546 42854
rect 484782 42618 484866 42854
rect 485102 42618 504546 42854
rect 504782 42618 504866 42854
rect 505102 42618 524546 42854
rect 524782 42618 524866 42854
rect 525102 42618 544546 42854
rect 544782 42618 544866 42854
rect 545102 42618 564546 42854
rect 564782 42618 564866 42854
rect 565102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 826 39454
rect 1062 39218 1146 39454
rect 1382 39218 24250 39454
rect 24486 39218 54970 39454
rect 55206 39218 80826 39454
rect 81062 39218 81146 39454
rect 81382 39218 100826 39454
rect 101062 39218 101146 39454
rect 101382 39218 120826 39454
rect 121062 39218 121146 39454
rect 121382 39218 140826 39454
rect 141062 39218 141146 39454
rect 141382 39218 160826 39454
rect 161062 39218 161146 39454
rect 161382 39218 180826 39454
rect 181062 39218 181146 39454
rect 181382 39218 200826 39454
rect 201062 39218 201146 39454
rect 201382 39218 220826 39454
rect 221062 39218 221146 39454
rect 221382 39218 240826 39454
rect 241062 39218 241146 39454
rect 241382 39218 260826 39454
rect 261062 39218 261146 39454
rect 261382 39218 280826 39454
rect 281062 39218 281146 39454
rect 281382 39218 300826 39454
rect 301062 39218 301146 39454
rect 301382 39218 320826 39454
rect 321062 39218 321146 39454
rect 321382 39218 340826 39454
rect 341062 39218 341146 39454
rect 341382 39218 360826 39454
rect 361062 39218 361146 39454
rect 361382 39218 380826 39454
rect 381062 39218 381146 39454
rect 381382 39218 400826 39454
rect 401062 39218 401146 39454
rect 401382 39218 420826 39454
rect 421062 39218 421146 39454
rect 421382 39218 440826 39454
rect 441062 39218 441146 39454
rect 441382 39218 460826 39454
rect 461062 39218 461146 39454
rect 461382 39218 480826 39454
rect 481062 39218 481146 39454
rect 481382 39218 500826 39454
rect 501062 39218 501146 39454
rect 501382 39218 520826 39454
rect 521062 39218 521146 39454
rect 521382 39218 540826 39454
rect 541062 39218 541146 39454
rect 541382 39218 560826 39454
rect 561062 39218 561146 39454
rect 561382 39218 580826 39454
rect 581062 39218 581146 39454
rect 581382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 826 39134
rect 1062 38898 1146 39134
rect 1382 38898 24250 39134
rect 24486 38898 54970 39134
rect 55206 38898 80826 39134
rect 81062 38898 81146 39134
rect 81382 38898 100826 39134
rect 101062 38898 101146 39134
rect 101382 38898 120826 39134
rect 121062 38898 121146 39134
rect 121382 38898 140826 39134
rect 141062 38898 141146 39134
rect 141382 38898 160826 39134
rect 161062 38898 161146 39134
rect 161382 38898 180826 39134
rect 181062 38898 181146 39134
rect 181382 38898 200826 39134
rect 201062 38898 201146 39134
rect 201382 38898 220826 39134
rect 221062 38898 221146 39134
rect 221382 38898 240826 39134
rect 241062 38898 241146 39134
rect 241382 38898 260826 39134
rect 261062 38898 261146 39134
rect 261382 38898 280826 39134
rect 281062 38898 281146 39134
rect 281382 38898 300826 39134
rect 301062 38898 301146 39134
rect 301382 38898 320826 39134
rect 321062 38898 321146 39134
rect 321382 38898 340826 39134
rect 341062 38898 341146 39134
rect 341382 38898 360826 39134
rect 361062 38898 361146 39134
rect 361382 38898 380826 39134
rect 381062 38898 381146 39134
rect 381382 38898 400826 39134
rect 401062 38898 401146 39134
rect 401382 38898 420826 39134
rect 421062 38898 421146 39134
rect 421382 38898 440826 39134
rect 441062 38898 441146 39134
rect 441382 38898 460826 39134
rect 461062 38898 461146 39134
rect 461382 38898 480826 39134
rect 481062 38898 481146 39134
rect 481382 38898 500826 39134
rect 501062 38898 501146 39134
rect 501382 38898 520826 39134
rect 521062 38898 521146 39134
rect 521382 38898 540826 39134
rect 541062 38898 541146 39134
rect 541382 38898 560826 39134
rect 561062 38898 561146 39134
rect 561382 38898 580826 39134
rect 581062 38898 581146 39134
rect 581382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 81986 32614
rect 82222 32378 82306 32614
rect 82542 32378 101986 32614
rect 102222 32378 102306 32614
rect 102542 32378 121986 32614
rect 122222 32378 122306 32614
rect 122542 32378 141986 32614
rect 142222 32378 142306 32614
rect 142542 32378 161986 32614
rect 162222 32378 162306 32614
rect 162542 32378 181986 32614
rect 182222 32378 182306 32614
rect 182542 32378 201986 32614
rect 202222 32378 202306 32614
rect 202542 32378 221986 32614
rect 222222 32378 222306 32614
rect 222542 32378 241986 32614
rect 242222 32378 242306 32614
rect 242542 32378 261986 32614
rect 262222 32378 262306 32614
rect 262542 32378 281986 32614
rect 282222 32378 282306 32614
rect 282542 32378 301986 32614
rect 302222 32378 302306 32614
rect 302542 32378 321986 32614
rect 322222 32378 322306 32614
rect 322542 32378 341986 32614
rect 342222 32378 342306 32614
rect 342542 32378 361986 32614
rect 362222 32378 362306 32614
rect 362542 32378 381986 32614
rect 382222 32378 382306 32614
rect 382542 32378 401986 32614
rect 402222 32378 402306 32614
rect 402542 32378 421986 32614
rect 422222 32378 422306 32614
rect 422542 32378 441986 32614
rect 442222 32378 442306 32614
rect 442542 32378 461986 32614
rect 462222 32378 462306 32614
rect 462542 32378 481986 32614
rect 482222 32378 482306 32614
rect 482542 32378 501986 32614
rect 502222 32378 502306 32614
rect 502542 32378 521986 32614
rect 522222 32378 522306 32614
rect 522542 32378 541986 32614
rect 542222 32378 542306 32614
rect 542542 32378 561986 32614
rect 562222 32378 562306 32614
rect 562542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 81986 32294
rect 82222 32058 82306 32294
rect 82542 32058 101986 32294
rect 102222 32058 102306 32294
rect 102542 32058 121986 32294
rect 122222 32058 122306 32294
rect 122542 32058 141986 32294
rect 142222 32058 142306 32294
rect 142542 32058 161986 32294
rect 162222 32058 162306 32294
rect 162542 32058 181986 32294
rect 182222 32058 182306 32294
rect 182542 32058 201986 32294
rect 202222 32058 202306 32294
rect 202542 32058 221986 32294
rect 222222 32058 222306 32294
rect 222542 32058 241986 32294
rect 242222 32058 242306 32294
rect 242542 32058 261986 32294
rect 262222 32058 262306 32294
rect 262542 32058 281986 32294
rect 282222 32058 282306 32294
rect 282542 32058 301986 32294
rect 302222 32058 302306 32294
rect 302542 32058 321986 32294
rect 322222 32058 322306 32294
rect 322542 32058 341986 32294
rect 342222 32058 342306 32294
rect 342542 32058 361986 32294
rect 362222 32058 362306 32294
rect 362542 32058 381986 32294
rect 382222 32058 382306 32294
rect 382542 32058 401986 32294
rect 402222 32058 402306 32294
rect 402542 32058 421986 32294
rect 422222 32058 422306 32294
rect 422542 32058 441986 32294
rect 442222 32058 442306 32294
rect 442542 32058 461986 32294
rect 462222 32058 462306 32294
rect 462542 32058 481986 32294
rect 482222 32058 482306 32294
rect 482542 32058 501986 32294
rect 502222 32058 502306 32294
rect 502542 32058 521986 32294
rect 522222 32058 522306 32294
rect 522542 32058 541986 32294
rect 542222 32058 542306 32294
rect 542542 32058 561986 32294
rect 562222 32058 562306 32294
rect 562542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 78266 28894
rect 78502 28658 78586 28894
rect 78822 28658 98266 28894
rect 98502 28658 98586 28894
rect 98822 28658 118266 28894
rect 118502 28658 118586 28894
rect 118822 28658 138266 28894
rect 138502 28658 138586 28894
rect 138822 28658 158266 28894
rect 158502 28658 158586 28894
rect 158822 28658 178266 28894
rect 178502 28658 178586 28894
rect 178822 28658 198266 28894
rect 198502 28658 198586 28894
rect 198822 28658 218266 28894
rect 218502 28658 218586 28894
rect 218822 28658 238266 28894
rect 238502 28658 238586 28894
rect 238822 28658 258266 28894
rect 258502 28658 258586 28894
rect 258822 28658 278266 28894
rect 278502 28658 278586 28894
rect 278822 28658 298266 28894
rect 298502 28658 298586 28894
rect 298822 28658 318266 28894
rect 318502 28658 318586 28894
rect 318822 28658 338266 28894
rect 338502 28658 338586 28894
rect 338822 28658 358266 28894
rect 358502 28658 358586 28894
rect 358822 28658 378266 28894
rect 378502 28658 378586 28894
rect 378822 28658 398266 28894
rect 398502 28658 398586 28894
rect 398822 28658 418266 28894
rect 418502 28658 418586 28894
rect 418822 28658 438266 28894
rect 438502 28658 438586 28894
rect 438822 28658 458266 28894
rect 458502 28658 458586 28894
rect 458822 28658 478266 28894
rect 478502 28658 478586 28894
rect 478822 28658 498266 28894
rect 498502 28658 498586 28894
rect 498822 28658 518266 28894
rect 518502 28658 518586 28894
rect 518822 28658 538266 28894
rect 538502 28658 538586 28894
rect 538822 28658 558266 28894
rect 558502 28658 558586 28894
rect 558822 28658 578266 28894
rect 578502 28658 578586 28894
rect 578822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 78266 28574
rect 78502 28338 78586 28574
rect 78822 28338 98266 28574
rect 98502 28338 98586 28574
rect 98822 28338 118266 28574
rect 118502 28338 118586 28574
rect 118822 28338 138266 28574
rect 138502 28338 138586 28574
rect 138822 28338 158266 28574
rect 158502 28338 158586 28574
rect 158822 28338 178266 28574
rect 178502 28338 178586 28574
rect 178822 28338 198266 28574
rect 198502 28338 198586 28574
rect 198822 28338 218266 28574
rect 218502 28338 218586 28574
rect 218822 28338 238266 28574
rect 238502 28338 238586 28574
rect 238822 28338 258266 28574
rect 258502 28338 258586 28574
rect 258822 28338 278266 28574
rect 278502 28338 278586 28574
rect 278822 28338 298266 28574
rect 298502 28338 298586 28574
rect 298822 28338 318266 28574
rect 318502 28338 318586 28574
rect 318822 28338 338266 28574
rect 338502 28338 338586 28574
rect 338822 28338 358266 28574
rect 358502 28338 358586 28574
rect 358822 28338 378266 28574
rect 378502 28338 378586 28574
rect 378822 28338 398266 28574
rect 398502 28338 398586 28574
rect 398822 28338 418266 28574
rect 418502 28338 418586 28574
rect 418822 28338 438266 28574
rect 438502 28338 438586 28574
rect 438822 28338 458266 28574
rect 458502 28338 458586 28574
rect 458822 28338 478266 28574
rect 478502 28338 478586 28574
rect 478822 28338 498266 28574
rect 498502 28338 498586 28574
rect 498822 28338 518266 28574
rect 518502 28338 518586 28574
rect 518822 28338 538266 28574
rect 538502 28338 538586 28574
rect 538822 28338 558266 28574
rect 558502 28338 558586 28574
rect 558822 28338 578266 28574
rect 578502 28338 578586 28574
rect 578822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 14546 25174
rect 14782 24938 14866 25174
rect 15102 24938 74546 25174
rect 74782 24938 74866 25174
rect 75102 24938 94546 25174
rect 94782 24938 94866 25174
rect 95102 24938 114546 25174
rect 114782 24938 114866 25174
rect 115102 24938 134546 25174
rect 134782 24938 134866 25174
rect 135102 24938 154546 25174
rect 154782 24938 154866 25174
rect 155102 24938 174546 25174
rect 174782 24938 174866 25174
rect 175102 24938 194546 25174
rect 194782 24938 194866 25174
rect 195102 24938 214546 25174
rect 214782 24938 214866 25174
rect 215102 24938 234546 25174
rect 234782 24938 234866 25174
rect 235102 24938 254546 25174
rect 254782 24938 254866 25174
rect 255102 24938 274546 25174
rect 274782 24938 274866 25174
rect 275102 24938 294546 25174
rect 294782 24938 294866 25174
rect 295102 24938 314546 25174
rect 314782 24938 314866 25174
rect 315102 24938 334546 25174
rect 334782 24938 334866 25174
rect 335102 24938 354546 25174
rect 354782 24938 354866 25174
rect 355102 24938 374546 25174
rect 374782 24938 374866 25174
rect 375102 24938 394546 25174
rect 394782 24938 394866 25174
rect 395102 24938 414546 25174
rect 414782 24938 414866 25174
rect 415102 24938 434546 25174
rect 434782 24938 434866 25174
rect 435102 24938 454546 25174
rect 454782 24938 454866 25174
rect 455102 24938 474546 25174
rect 474782 24938 474866 25174
rect 475102 24938 494546 25174
rect 494782 24938 494866 25174
rect 495102 24938 514546 25174
rect 514782 24938 514866 25174
rect 515102 24938 534546 25174
rect 534782 24938 534866 25174
rect 535102 24938 554546 25174
rect 554782 24938 554866 25174
rect 555102 24938 574546 25174
rect 574782 24938 574866 25174
rect 575102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 14546 24854
rect 14782 24618 14866 24854
rect 15102 24618 74546 24854
rect 74782 24618 74866 24854
rect 75102 24618 94546 24854
rect 94782 24618 94866 24854
rect 95102 24618 114546 24854
rect 114782 24618 114866 24854
rect 115102 24618 134546 24854
rect 134782 24618 134866 24854
rect 135102 24618 154546 24854
rect 154782 24618 154866 24854
rect 155102 24618 174546 24854
rect 174782 24618 174866 24854
rect 175102 24618 194546 24854
rect 194782 24618 194866 24854
rect 195102 24618 214546 24854
rect 214782 24618 214866 24854
rect 215102 24618 234546 24854
rect 234782 24618 234866 24854
rect 235102 24618 254546 24854
rect 254782 24618 254866 24854
rect 255102 24618 274546 24854
rect 274782 24618 274866 24854
rect 275102 24618 294546 24854
rect 294782 24618 294866 24854
rect 295102 24618 314546 24854
rect 314782 24618 314866 24854
rect 315102 24618 334546 24854
rect 334782 24618 334866 24854
rect 335102 24618 354546 24854
rect 354782 24618 354866 24854
rect 355102 24618 374546 24854
rect 374782 24618 374866 24854
rect 375102 24618 394546 24854
rect 394782 24618 394866 24854
rect 395102 24618 414546 24854
rect 414782 24618 414866 24854
rect 415102 24618 434546 24854
rect 434782 24618 434866 24854
rect 435102 24618 454546 24854
rect 454782 24618 454866 24854
rect 455102 24618 474546 24854
rect 474782 24618 474866 24854
rect 475102 24618 494546 24854
rect 494782 24618 494866 24854
rect 495102 24618 514546 24854
rect 514782 24618 514866 24854
rect 515102 24618 534546 24854
rect 534782 24618 534866 24854
rect 535102 24618 554546 24854
rect 554782 24618 554866 24854
rect 555102 24618 574546 24854
rect 574782 24618 574866 24854
rect 575102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 10826 21454
rect 11062 21218 11146 21454
rect 11382 21218 90826 21454
rect 91062 21218 91146 21454
rect 91382 21218 110826 21454
rect 111062 21218 111146 21454
rect 111382 21218 130826 21454
rect 131062 21218 131146 21454
rect 131382 21218 150826 21454
rect 151062 21218 151146 21454
rect 151382 21218 170826 21454
rect 171062 21218 171146 21454
rect 171382 21218 190826 21454
rect 191062 21218 191146 21454
rect 191382 21218 210826 21454
rect 211062 21218 211146 21454
rect 211382 21218 230826 21454
rect 231062 21218 231146 21454
rect 231382 21218 250826 21454
rect 251062 21218 251146 21454
rect 251382 21218 270826 21454
rect 271062 21218 271146 21454
rect 271382 21218 290826 21454
rect 291062 21218 291146 21454
rect 291382 21218 310826 21454
rect 311062 21218 311146 21454
rect 311382 21218 330826 21454
rect 331062 21218 331146 21454
rect 331382 21218 350826 21454
rect 351062 21218 351146 21454
rect 351382 21218 370826 21454
rect 371062 21218 371146 21454
rect 371382 21218 390826 21454
rect 391062 21218 391146 21454
rect 391382 21218 410826 21454
rect 411062 21218 411146 21454
rect 411382 21218 430826 21454
rect 431062 21218 431146 21454
rect 431382 21218 450826 21454
rect 451062 21218 451146 21454
rect 451382 21218 470826 21454
rect 471062 21218 471146 21454
rect 471382 21218 490826 21454
rect 491062 21218 491146 21454
rect 491382 21218 510826 21454
rect 511062 21218 511146 21454
rect 511382 21218 530826 21454
rect 531062 21218 531146 21454
rect 531382 21218 550826 21454
rect 551062 21218 551146 21454
rect 551382 21218 570826 21454
rect 571062 21218 571146 21454
rect 571382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 10826 21134
rect 11062 20898 11146 21134
rect 11382 20898 90826 21134
rect 91062 20898 91146 21134
rect 91382 20898 110826 21134
rect 111062 20898 111146 21134
rect 111382 20898 130826 21134
rect 131062 20898 131146 21134
rect 131382 20898 150826 21134
rect 151062 20898 151146 21134
rect 151382 20898 170826 21134
rect 171062 20898 171146 21134
rect 171382 20898 190826 21134
rect 191062 20898 191146 21134
rect 191382 20898 210826 21134
rect 211062 20898 211146 21134
rect 211382 20898 230826 21134
rect 231062 20898 231146 21134
rect 231382 20898 250826 21134
rect 251062 20898 251146 21134
rect 251382 20898 270826 21134
rect 271062 20898 271146 21134
rect 271382 20898 290826 21134
rect 291062 20898 291146 21134
rect 291382 20898 310826 21134
rect 311062 20898 311146 21134
rect 311382 20898 330826 21134
rect 331062 20898 331146 21134
rect 331382 20898 350826 21134
rect 351062 20898 351146 21134
rect 351382 20898 370826 21134
rect 371062 20898 371146 21134
rect 371382 20898 390826 21134
rect 391062 20898 391146 21134
rect 391382 20898 410826 21134
rect 411062 20898 411146 21134
rect 411382 20898 430826 21134
rect 431062 20898 431146 21134
rect 431382 20898 450826 21134
rect 451062 20898 451146 21134
rect 451382 20898 470826 21134
rect 471062 20898 471146 21134
rect 471382 20898 490826 21134
rect 491062 20898 491146 21134
rect 491382 20898 510826 21134
rect 511062 20898 511146 21134
rect 511382 20898 530826 21134
rect 531062 20898 531146 21134
rect 531382 20898 550826 21134
rect 551062 20898 551146 21134
rect 551382 20898 570826 21134
rect 571062 20898 571146 21134
rect 571382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 11986 14614
rect 12222 14378 12306 14614
rect 12542 14378 31986 14614
rect 32222 14378 32306 14614
rect 32542 14378 51986 14614
rect 52222 14378 52306 14614
rect 52542 14378 71986 14614
rect 72222 14378 72306 14614
rect 72542 14378 91986 14614
rect 92222 14378 92306 14614
rect 92542 14378 111986 14614
rect 112222 14378 112306 14614
rect 112542 14378 131986 14614
rect 132222 14378 132306 14614
rect 132542 14378 151986 14614
rect 152222 14378 152306 14614
rect 152542 14378 171986 14614
rect 172222 14378 172306 14614
rect 172542 14378 191986 14614
rect 192222 14378 192306 14614
rect 192542 14378 211986 14614
rect 212222 14378 212306 14614
rect 212542 14378 231986 14614
rect 232222 14378 232306 14614
rect 232542 14378 251986 14614
rect 252222 14378 252306 14614
rect 252542 14378 271986 14614
rect 272222 14378 272306 14614
rect 272542 14378 291986 14614
rect 292222 14378 292306 14614
rect 292542 14378 311986 14614
rect 312222 14378 312306 14614
rect 312542 14378 331986 14614
rect 332222 14378 332306 14614
rect 332542 14378 351986 14614
rect 352222 14378 352306 14614
rect 352542 14378 371986 14614
rect 372222 14378 372306 14614
rect 372542 14378 391986 14614
rect 392222 14378 392306 14614
rect 392542 14378 411986 14614
rect 412222 14378 412306 14614
rect 412542 14378 431986 14614
rect 432222 14378 432306 14614
rect 432542 14378 451986 14614
rect 452222 14378 452306 14614
rect 452542 14378 471986 14614
rect 472222 14378 472306 14614
rect 472542 14378 491986 14614
rect 492222 14378 492306 14614
rect 492542 14378 511986 14614
rect 512222 14378 512306 14614
rect 512542 14378 531986 14614
rect 532222 14378 532306 14614
rect 532542 14378 551986 14614
rect 552222 14378 552306 14614
rect 552542 14378 571986 14614
rect 572222 14378 572306 14614
rect 572542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 11986 14294
rect 12222 14058 12306 14294
rect 12542 14058 31986 14294
rect 32222 14058 32306 14294
rect 32542 14058 51986 14294
rect 52222 14058 52306 14294
rect 52542 14058 71986 14294
rect 72222 14058 72306 14294
rect 72542 14058 91986 14294
rect 92222 14058 92306 14294
rect 92542 14058 111986 14294
rect 112222 14058 112306 14294
rect 112542 14058 131986 14294
rect 132222 14058 132306 14294
rect 132542 14058 151986 14294
rect 152222 14058 152306 14294
rect 152542 14058 171986 14294
rect 172222 14058 172306 14294
rect 172542 14058 191986 14294
rect 192222 14058 192306 14294
rect 192542 14058 211986 14294
rect 212222 14058 212306 14294
rect 212542 14058 231986 14294
rect 232222 14058 232306 14294
rect 232542 14058 251986 14294
rect 252222 14058 252306 14294
rect 252542 14058 271986 14294
rect 272222 14058 272306 14294
rect 272542 14058 291986 14294
rect 292222 14058 292306 14294
rect 292542 14058 311986 14294
rect 312222 14058 312306 14294
rect 312542 14058 331986 14294
rect 332222 14058 332306 14294
rect 332542 14058 351986 14294
rect 352222 14058 352306 14294
rect 352542 14058 371986 14294
rect 372222 14058 372306 14294
rect 372542 14058 391986 14294
rect 392222 14058 392306 14294
rect 392542 14058 411986 14294
rect 412222 14058 412306 14294
rect 412542 14058 431986 14294
rect 432222 14058 432306 14294
rect 432542 14058 451986 14294
rect 452222 14058 452306 14294
rect 452542 14058 471986 14294
rect 472222 14058 472306 14294
rect 472542 14058 491986 14294
rect 492222 14058 492306 14294
rect 492542 14058 511986 14294
rect 512222 14058 512306 14294
rect 512542 14058 531986 14294
rect 532222 14058 532306 14294
rect 532542 14058 551986 14294
rect 552222 14058 552306 14294
rect 552542 14058 571986 14294
rect 572222 14058 572306 14294
rect 572542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 8266 10894
rect 8502 10658 8586 10894
rect 8822 10658 28266 10894
rect 28502 10658 28586 10894
rect 28822 10658 48266 10894
rect 48502 10658 48586 10894
rect 48822 10658 68266 10894
rect 68502 10658 68586 10894
rect 68822 10658 88266 10894
rect 88502 10658 88586 10894
rect 88822 10658 108266 10894
rect 108502 10658 108586 10894
rect 108822 10658 128266 10894
rect 128502 10658 128586 10894
rect 128822 10658 148266 10894
rect 148502 10658 148586 10894
rect 148822 10658 168266 10894
rect 168502 10658 168586 10894
rect 168822 10658 188266 10894
rect 188502 10658 188586 10894
rect 188822 10658 208266 10894
rect 208502 10658 208586 10894
rect 208822 10658 228266 10894
rect 228502 10658 228586 10894
rect 228822 10658 248266 10894
rect 248502 10658 248586 10894
rect 248822 10658 268266 10894
rect 268502 10658 268586 10894
rect 268822 10658 288266 10894
rect 288502 10658 288586 10894
rect 288822 10658 308266 10894
rect 308502 10658 308586 10894
rect 308822 10658 328266 10894
rect 328502 10658 328586 10894
rect 328822 10658 348266 10894
rect 348502 10658 348586 10894
rect 348822 10658 368266 10894
rect 368502 10658 368586 10894
rect 368822 10658 388266 10894
rect 388502 10658 388586 10894
rect 388822 10658 408266 10894
rect 408502 10658 408586 10894
rect 408822 10658 428266 10894
rect 428502 10658 428586 10894
rect 428822 10658 448266 10894
rect 448502 10658 448586 10894
rect 448822 10658 468266 10894
rect 468502 10658 468586 10894
rect 468822 10658 488266 10894
rect 488502 10658 488586 10894
rect 488822 10658 508266 10894
rect 508502 10658 508586 10894
rect 508822 10658 528266 10894
rect 528502 10658 528586 10894
rect 528822 10658 548266 10894
rect 548502 10658 548586 10894
rect 548822 10658 568266 10894
rect 568502 10658 568586 10894
rect 568822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 8266 10574
rect 8502 10338 8586 10574
rect 8822 10338 28266 10574
rect 28502 10338 28586 10574
rect 28822 10338 48266 10574
rect 48502 10338 48586 10574
rect 48822 10338 68266 10574
rect 68502 10338 68586 10574
rect 68822 10338 88266 10574
rect 88502 10338 88586 10574
rect 88822 10338 108266 10574
rect 108502 10338 108586 10574
rect 108822 10338 128266 10574
rect 128502 10338 128586 10574
rect 128822 10338 148266 10574
rect 148502 10338 148586 10574
rect 148822 10338 168266 10574
rect 168502 10338 168586 10574
rect 168822 10338 188266 10574
rect 188502 10338 188586 10574
rect 188822 10338 208266 10574
rect 208502 10338 208586 10574
rect 208822 10338 228266 10574
rect 228502 10338 228586 10574
rect 228822 10338 248266 10574
rect 248502 10338 248586 10574
rect 248822 10338 268266 10574
rect 268502 10338 268586 10574
rect 268822 10338 288266 10574
rect 288502 10338 288586 10574
rect 288822 10338 308266 10574
rect 308502 10338 308586 10574
rect 308822 10338 328266 10574
rect 328502 10338 328586 10574
rect 328822 10338 348266 10574
rect 348502 10338 348586 10574
rect 348822 10338 368266 10574
rect 368502 10338 368586 10574
rect 368822 10338 388266 10574
rect 388502 10338 388586 10574
rect 388822 10338 408266 10574
rect 408502 10338 408586 10574
rect 408822 10338 428266 10574
rect 428502 10338 428586 10574
rect 428822 10338 448266 10574
rect 448502 10338 448586 10574
rect 448822 10338 468266 10574
rect 468502 10338 468586 10574
rect 468822 10338 488266 10574
rect 488502 10338 488586 10574
rect 488822 10338 508266 10574
rect 508502 10338 508586 10574
rect 508822 10338 528266 10574
rect 528502 10338 528586 10574
rect 528822 10338 548266 10574
rect 548502 10338 548586 10574
rect 548822 10338 568266 10574
rect 568502 10338 568586 10574
rect 568822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 4546 7174
rect 4782 6938 4866 7174
rect 5102 6938 24546 7174
rect 24782 6938 24866 7174
rect 25102 6938 44546 7174
rect 44782 6938 44866 7174
rect 45102 6938 64546 7174
rect 64782 6938 64866 7174
rect 65102 6938 84546 7174
rect 84782 6938 84866 7174
rect 85102 6938 104546 7174
rect 104782 6938 104866 7174
rect 105102 6938 124546 7174
rect 124782 6938 124866 7174
rect 125102 6938 144546 7174
rect 144782 6938 144866 7174
rect 145102 6938 164546 7174
rect 164782 6938 164866 7174
rect 165102 6938 184546 7174
rect 184782 6938 184866 7174
rect 185102 6938 204546 7174
rect 204782 6938 204866 7174
rect 205102 6938 224546 7174
rect 224782 6938 224866 7174
rect 225102 6938 244546 7174
rect 244782 6938 244866 7174
rect 245102 6938 264546 7174
rect 264782 6938 264866 7174
rect 265102 6938 284546 7174
rect 284782 6938 284866 7174
rect 285102 6938 304546 7174
rect 304782 6938 304866 7174
rect 305102 6938 324546 7174
rect 324782 6938 324866 7174
rect 325102 6938 344546 7174
rect 344782 6938 344866 7174
rect 345102 6938 364546 7174
rect 364782 6938 364866 7174
rect 365102 6938 384546 7174
rect 384782 6938 384866 7174
rect 385102 6938 404546 7174
rect 404782 6938 404866 7174
rect 405102 6938 424546 7174
rect 424782 6938 424866 7174
rect 425102 6938 444546 7174
rect 444782 6938 444866 7174
rect 445102 6938 464546 7174
rect 464782 6938 464866 7174
rect 465102 6938 484546 7174
rect 484782 6938 484866 7174
rect 485102 6938 504546 7174
rect 504782 6938 504866 7174
rect 505102 6938 524546 7174
rect 524782 6938 524866 7174
rect 525102 6938 544546 7174
rect 544782 6938 544866 7174
rect 545102 6938 564546 7174
rect 564782 6938 564866 7174
rect 565102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 4546 6854
rect 4782 6618 4866 6854
rect 5102 6618 24546 6854
rect 24782 6618 24866 6854
rect 25102 6618 44546 6854
rect 44782 6618 44866 6854
rect 45102 6618 64546 6854
rect 64782 6618 64866 6854
rect 65102 6618 84546 6854
rect 84782 6618 84866 6854
rect 85102 6618 104546 6854
rect 104782 6618 104866 6854
rect 105102 6618 124546 6854
rect 124782 6618 124866 6854
rect 125102 6618 144546 6854
rect 144782 6618 144866 6854
rect 145102 6618 164546 6854
rect 164782 6618 164866 6854
rect 165102 6618 184546 6854
rect 184782 6618 184866 6854
rect 185102 6618 204546 6854
rect 204782 6618 204866 6854
rect 205102 6618 224546 6854
rect 224782 6618 224866 6854
rect 225102 6618 244546 6854
rect 244782 6618 244866 6854
rect 245102 6618 264546 6854
rect 264782 6618 264866 6854
rect 265102 6618 284546 6854
rect 284782 6618 284866 6854
rect 285102 6618 304546 6854
rect 304782 6618 304866 6854
rect 305102 6618 324546 6854
rect 324782 6618 324866 6854
rect 325102 6618 344546 6854
rect 344782 6618 344866 6854
rect 345102 6618 364546 6854
rect 364782 6618 364866 6854
rect 365102 6618 384546 6854
rect 384782 6618 384866 6854
rect 385102 6618 404546 6854
rect 404782 6618 404866 6854
rect 405102 6618 424546 6854
rect 424782 6618 424866 6854
rect 425102 6618 444546 6854
rect 444782 6618 444866 6854
rect 445102 6618 464546 6854
rect 464782 6618 464866 6854
rect 465102 6618 484546 6854
rect 484782 6618 484866 6854
rect 485102 6618 504546 6854
rect 504782 6618 504866 6854
rect 505102 6618 524546 6854
rect 524782 6618 524866 6854
rect 525102 6618 544546 6854
rect 544782 6618 544866 6854
rect 545102 6618 564546 6854
rect 564782 6618 564866 6854
rect 565102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 826 3454
rect 1062 3218 1146 3454
rect 1382 3218 20826 3454
rect 21062 3218 21146 3454
rect 21382 3218 40826 3454
rect 41062 3218 41146 3454
rect 41382 3218 60826 3454
rect 61062 3218 61146 3454
rect 61382 3218 80826 3454
rect 81062 3218 81146 3454
rect 81382 3218 100826 3454
rect 101062 3218 101146 3454
rect 101382 3218 120826 3454
rect 121062 3218 121146 3454
rect 121382 3218 140826 3454
rect 141062 3218 141146 3454
rect 141382 3218 160826 3454
rect 161062 3218 161146 3454
rect 161382 3218 180826 3454
rect 181062 3218 181146 3454
rect 181382 3218 200826 3454
rect 201062 3218 201146 3454
rect 201382 3218 220826 3454
rect 221062 3218 221146 3454
rect 221382 3218 240826 3454
rect 241062 3218 241146 3454
rect 241382 3218 260826 3454
rect 261062 3218 261146 3454
rect 261382 3218 280826 3454
rect 281062 3218 281146 3454
rect 281382 3218 300826 3454
rect 301062 3218 301146 3454
rect 301382 3218 320826 3454
rect 321062 3218 321146 3454
rect 321382 3218 340826 3454
rect 341062 3218 341146 3454
rect 341382 3218 360826 3454
rect 361062 3218 361146 3454
rect 361382 3218 380826 3454
rect 381062 3218 381146 3454
rect 381382 3218 400826 3454
rect 401062 3218 401146 3454
rect 401382 3218 420826 3454
rect 421062 3218 421146 3454
rect 421382 3218 440826 3454
rect 441062 3218 441146 3454
rect 441382 3218 460826 3454
rect 461062 3218 461146 3454
rect 461382 3218 480826 3454
rect 481062 3218 481146 3454
rect 481382 3218 500826 3454
rect 501062 3218 501146 3454
rect 501382 3218 520826 3454
rect 521062 3218 521146 3454
rect 521382 3218 540826 3454
rect 541062 3218 541146 3454
rect 541382 3218 560826 3454
rect 561062 3218 561146 3454
rect 561382 3218 580826 3454
rect 581062 3218 581146 3454
rect 581382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 826 3134
rect 1062 2898 1146 3134
rect 1382 2898 20826 3134
rect 21062 2898 21146 3134
rect 21382 2898 40826 3134
rect 41062 2898 41146 3134
rect 41382 2898 60826 3134
rect 61062 2898 61146 3134
rect 61382 2898 80826 3134
rect 81062 2898 81146 3134
rect 81382 2898 100826 3134
rect 101062 2898 101146 3134
rect 101382 2898 120826 3134
rect 121062 2898 121146 3134
rect 121382 2898 140826 3134
rect 141062 2898 141146 3134
rect 141382 2898 160826 3134
rect 161062 2898 161146 3134
rect 161382 2898 180826 3134
rect 181062 2898 181146 3134
rect 181382 2898 200826 3134
rect 201062 2898 201146 3134
rect 201382 2898 220826 3134
rect 221062 2898 221146 3134
rect 221382 2898 240826 3134
rect 241062 2898 241146 3134
rect 241382 2898 260826 3134
rect 261062 2898 261146 3134
rect 261382 2898 280826 3134
rect 281062 2898 281146 3134
rect 281382 2898 300826 3134
rect 301062 2898 301146 3134
rect 301382 2898 320826 3134
rect 321062 2898 321146 3134
rect 321382 2898 340826 3134
rect 341062 2898 341146 3134
rect 341382 2898 360826 3134
rect 361062 2898 361146 3134
rect 361382 2898 380826 3134
rect 381062 2898 381146 3134
rect 381382 2898 400826 3134
rect 401062 2898 401146 3134
rect 401382 2898 420826 3134
rect 421062 2898 421146 3134
rect 421382 2898 440826 3134
rect 441062 2898 441146 3134
rect 441382 2898 460826 3134
rect 461062 2898 461146 3134
rect 461382 2898 480826 3134
rect 481062 2898 481146 3134
rect 481382 2898 500826 3134
rect 501062 2898 501146 3134
rect 501382 2898 520826 3134
rect 521062 2898 521146 3134
rect 521382 2898 540826 3134
rect 541062 2898 541146 3134
rect 541382 2898 560826 3134
rect 561062 2898 561146 3134
rect 561382 2898 580826 3134
rect 581062 2898 581146 3134
rect 581382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 826 -346
rect 1062 -582 1146 -346
rect 1382 -582 20826 -346
rect 21062 -582 21146 -346
rect 21382 -582 40826 -346
rect 41062 -582 41146 -346
rect 41382 -582 60826 -346
rect 61062 -582 61146 -346
rect 61382 -582 80826 -346
rect 81062 -582 81146 -346
rect 81382 -582 100826 -346
rect 101062 -582 101146 -346
rect 101382 -582 120826 -346
rect 121062 -582 121146 -346
rect 121382 -582 140826 -346
rect 141062 -582 141146 -346
rect 141382 -582 160826 -346
rect 161062 -582 161146 -346
rect 161382 -582 180826 -346
rect 181062 -582 181146 -346
rect 181382 -582 200826 -346
rect 201062 -582 201146 -346
rect 201382 -582 220826 -346
rect 221062 -582 221146 -346
rect 221382 -582 240826 -346
rect 241062 -582 241146 -346
rect 241382 -582 260826 -346
rect 261062 -582 261146 -346
rect 261382 -582 280826 -346
rect 281062 -582 281146 -346
rect 281382 -582 300826 -346
rect 301062 -582 301146 -346
rect 301382 -582 320826 -346
rect 321062 -582 321146 -346
rect 321382 -582 340826 -346
rect 341062 -582 341146 -346
rect 341382 -582 360826 -346
rect 361062 -582 361146 -346
rect 361382 -582 380826 -346
rect 381062 -582 381146 -346
rect 381382 -582 400826 -346
rect 401062 -582 401146 -346
rect 401382 -582 420826 -346
rect 421062 -582 421146 -346
rect 421382 -582 440826 -346
rect 441062 -582 441146 -346
rect 441382 -582 460826 -346
rect 461062 -582 461146 -346
rect 461382 -582 480826 -346
rect 481062 -582 481146 -346
rect 481382 -582 500826 -346
rect 501062 -582 501146 -346
rect 501382 -582 520826 -346
rect 521062 -582 521146 -346
rect 521382 -582 540826 -346
rect 541062 -582 541146 -346
rect 541382 -582 560826 -346
rect 561062 -582 561146 -346
rect 561382 -582 580826 -346
rect 581062 -582 581146 -346
rect 581382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 826 -666
rect 1062 -902 1146 -666
rect 1382 -902 20826 -666
rect 21062 -902 21146 -666
rect 21382 -902 40826 -666
rect 41062 -902 41146 -666
rect 41382 -902 60826 -666
rect 61062 -902 61146 -666
rect 61382 -902 80826 -666
rect 81062 -902 81146 -666
rect 81382 -902 100826 -666
rect 101062 -902 101146 -666
rect 101382 -902 120826 -666
rect 121062 -902 121146 -666
rect 121382 -902 140826 -666
rect 141062 -902 141146 -666
rect 141382 -902 160826 -666
rect 161062 -902 161146 -666
rect 161382 -902 180826 -666
rect 181062 -902 181146 -666
rect 181382 -902 200826 -666
rect 201062 -902 201146 -666
rect 201382 -902 220826 -666
rect 221062 -902 221146 -666
rect 221382 -902 240826 -666
rect 241062 -902 241146 -666
rect 241382 -902 260826 -666
rect 261062 -902 261146 -666
rect 261382 -902 280826 -666
rect 281062 -902 281146 -666
rect 281382 -902 300826 -666
rect 301062 -902 301146 -666
rect 301382 -902 320826 -666
rect 321062 -902 321146 -666
rect 321382 -902 340826 -666
rect 341062 -902 341146 -666
rect 341382 -902 360826 -666
rect 361062 -902 361146 -666
rect 361382 -902 380826 -666
rect 381062 -902 381146 -666
rect 381382 -902 400826 -666
rect 401062 -902 401146 -666
rect 401382 -902 420826 -666
rect 421062 -902 421146 -666
rect 421382 -902 440826 -666
rect 441062 -902 441146 -666
rect 441382 -902 460826 -666
rect 461062 -902 461146 -666
rect 461382 -902 480826 -666
rect 481062 -902 481146 -666
rect 481382 -902 500826 -666
rect 501062 -902 501146 -666
rect 501382 -902 520826 -666
rect 521062 -902 521146 -666
rect 521382 -902 540826 -666
rect 541062 -902 541146 -666
rect 541382 -902 560826 -666
rect 561062 -902 561146 -666
rect 561382 -902 580826 -666
rect 581062 -902 581146 -666
rect 581382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 10826 -1306
rect 11062 -1542 11146 -1306
rect 11382 -1542 30826 -1306
rect 31062 -1542 31146 -1306
rect 31382 -1542 50826 -1306
rect 51062 -1542 51146 -1306
rect 51382 -1542 70826 -1306
rect 71062 -1542 71146 -1306
rect 71382 -1542 90826 -1306
rect 91062 -1542 91146 -1306
rect 91382 -1542 110826 -1306
rect 111062 -1542 111146 -1306
rect 111382 -1542 130826 -1306
rect 131062 -1542 131146 -1306
rect 131382 -1542 150826 -1306
rect 151062 -1542 151146 -1306
rect 151382 -1542 170826 -1306
rect 171062 -1542 171146 -1306
rect 171382 -1542 190826 -1306
rect 191062 -1542 191146 -1306
rect 191382 -1542 210826 -1306
rect 211062 -1542 211146 -1306
rect 211382 -1542 230826 -1306
rect 231062 -1542 231146 -1306
rect 231382 -1542 250826 -1306
rect 251062 -1542 251146 -1306
rect 251382 -1542 270826 -1306
rect 271062 -1542 271146 -1306
rect 271382 -1542 290826 -1306
rect 291062 -1542 291146 -1306
rect 291382 -1542 310826 -1306
rect 311062 -1542 311146 -1306
rect 311382 -1542 330826 -1306
rect 331062 -1542 331146 -1306
rect 331382 -1542 350826 -1306
rect 351062 -1542 351146 -1306
rect 351382 -1542 370826 -1306
rect 371062 -1542 371146 -1306
rect 371382 -1542 390826 -1306
rect 391062 -1542 391146 -1306
rect 391382 -1542 410826 -1306
rect 411062 -1542 411146 -1306
rect 411382 -1542 430826 -1306
rect 431062 -1542 431146 -1306
rect 431382 -1542 450826 -1306
rect 451062 -1542 451146 -1306
rect 451382 -1542 470826 -1306
rect 471062 -1542 471146 -1306
rect 471382 -1542 490826 -1306
rect 491062 -1542 491146 -1306
rect 491382 -1542 510826 -1306
rect 511062 -1542 511146 -1306
rect 511382 -1542 530826 -1306
rect 531062 -1542 531146 -1306
rect 531382 -1542 550826 -1306
rect 551062 -1542 551146 -1306
rect 551382 -1542 570826 -1306
rect 571062 -1542 571146 -1306
rect 571382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 10826 -1626
rect 11062 -1862 11146 -1626
rect 11382 -1862 30826 -1626
rect 31062 -1862 31146 -1626
rect 31382 -1862 50826 -1626
rect 51062 -1862 51146 -1626
rect 51382 -1862 70826 -1626
rect 71062 -1862 71146 -1626
rect 71382 -1862 90826 -1626
rect 91062 -1862 91146 -1626
rect 91382 -1862 110826 -1626
rect 111062 -1862 111146 -1626
rect 111382 -1862 130826 -1626
rect 131062 -1862 131146 -1626
rect 131382 -1862 150826 -1626
rect 151062 -1862 151146 -1626
rect 151382 -1862 170826 -1626
rect 171062 -1862 171146 -1626
rect 171382 -1862 190826 -1626
rect 191062 -1862 191146 -1626
rect 191382 -1862 210826 -1626
rect 211062 -1862 211146 -1626
rect 211382 -1862 230826 -1626
rect 231062 -1862 231146 -1626
rect 231382 -1862 250826 -1626
rect 251062 -1862 251146 -1626
rect 251382 -1862 270826 -1626
rect 271062 -1862 271146 -1626
rect 271382 -1862 290826 -1626
rect 291062 -1862 291146 -1626
rect 291382 -1862 310826 -1626
rect 311062 -1862 311146 -1626
rect 311382 -1862 330826 -1626
rect 331062 -1862 331146 -1626
rect 331382 -1862 350826 -1626
rect 351062 -1862 351146 -1626
rect 351382 -1862 370826 -1626
rect 371062 -1862 371146 -1626
rect 371382 -1862 390826 -1626
rect 391062 -1862 391146 -1626
rect 391382 -1862 410826 -1626
rect 411062 -1862 411146 -1626
rect 411382 -1862 430826 -1626
rect 431062 -1862 431146 -1626
rect 431382 -1862 450826 -1626
rect 451062 -1862 451146 -1626
rect 451382 -1862 470826 -1626
rect 471062 -1862 471146 -1626
rect 471382 -1862 490826 -1626
rect 491062 -1862 491146 -1626
rect 491382 -1862 510826 -1626
rect 511062 -1862 511146 -1626
rect 511382 -1862 530826 -1626
rect 531062 -1862 531146 -1626
rect 531382 -1862 550826 -1626
rect 551062 -1862 551146 -1626
rect 551382 -1862 570826 -1626
rect 571062 -1862 571146 -1626
rect 571382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 4546 -2266
rect 4782 -2502 4866 -2266
rect 5102 -2502 24546 -2266
rect 24782 -2502 24866 -2266
rect 25102 -2502 44546 -2266
rect 44782 -2502 44866 -2266
rect 45102 -2502 64546 -2266
rect 64782 -2502 64866 -2266
rect 65102 -2502 84546 -2266
rect 84782 -2502 84866 -2266
rect 85102 -2502 104546 -2266
rect 104782 -2502 104866 -2266
rect 105102 -2502 124546 -2266
rect 124782 -2502 124866 -2266
rect 125102 -2502 144546 -2266
rect 144782 -2502 144866 -2266
rect 145102 -2502 164546 -2266
rect 164782 -2502 164866 -2266
rect 165102 -2502 184546 -2266
rect 184782 -2502 184866 -2266
rect 185102 -2502 204546 -2266
rect 204782 -2502 204866 -2266
rect 205102 -2502 224546 -2266
rect 224782 -2502 224866 -2266
rect 225102 -2502 244546 -2266
rect 244782 -2502 244866 -2266
rect 245102 -2502 264546 -2266
rect 264782 -2502 264866 -2266
rect 265102 -2502 284546 -2266
rect 284782 -2502 284866 -2266
rect 285102 -2502 304546 -2266
rect 304782 -2502 304866 -2266
rect 305102 -2502 324546 -2266
rect 324782 -2502 324866 -2266
rect 325102 -2502 344546 -2266
rect 344782 -2502 344866 -2266
rect 345102 -2502 364546 -2266
rect 364782 -2502 364866 -2266
rect 365102 -2502 384546 -2266
rect 384782 -2502 384866 -2266
rect 385102 -2502 404546 -2266
rect 404782 -2502 404866 -2266
rect 405102 -2502 424546 -2266
rect 424782 -2502 424866 -2266
rect 425102 -2502 444546 -2266
rect 444782 -2502 444866 -2266
rect 445102 -2502 464546 -2266
rect 464782 -2502 464866 -2266
rect 465102 -2502 484546 -2266
rect 484782 -2502 484866 -2266
rect 485102 -2502 504546 -2266
rect 504782 -2502 504866 -2266
rect 505102 -2502 524546 -2266
rect 524782 -2502 524866 -2266
rect 525102 -2502 544546 -2266
rect 544782 -2502 544866 -2266
rect 545102 -2502 564546 -2266
rect 564782 -2502 564866 -2266
rect 565102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 4546 -2586
rect 4782 -2822 4866 -2586
rect 5102 -2822 24546 -2586
rect 24782 -2822 24866 -2586
rect 25102 -2822 44546 -2586
rect 44782 -2822 44866 -2586
rect 45102 -2822 64546 -2586
rect 64782 -2822 64866 -2586
rect 65102 -2822 84546 -2586
rect 84782 -2822 84866 -2586
rect 85102 -2822 104546 -2586
rect 104782 -2822 104866 -2586
rect 105102 -2822 124546 -2586
rect 124782 -2822 124866 -2586
rect 125102 -2822 144546 -2586
rect 144782 -2822 144866 -2586
rect 145102 -2822 164546 -2586
rect 164782 -2822 164866 -2586
rect 165102 -2822 184546 -2586
rect 184782 -2822 184866 -2586
rect 185102 -2822 204546 -2586
rect 204782 -2822 204866 -2586
rect 205102 -2822 224546 -2586
rect 224782 -2822 224866 -2586
rect 225102 -2822 244546 -2586
rect 244782 -2822 244866 -2586
rect 245102 -2822 264546 -2586
rect 264782 -2822 264866 -2586
rect 265102 -2822 284546 -2586
rect 284782 -2822 284866 -2586
rect 285102 -2822 304546 -2586
rect 304782 -2822 304866 -2586
rect 305102 -2822 324546 -2586
rect 324782 -2822 324866 -2586
rect 325102 -2822 344546 -2586
rect 344782 -2822 344866 -2586
rect 345102 -2822 364546 -2586
rect 364782 -2822 364866 -2586
rect 365102 -2822 384546 -2586
rect 384782 -2822 384866 -2586
rect 385102 -2822 404546 -2586
rect 404782 -2822 404866 -2586
rect 405102 -2822 424546 -2586
rect 424782 -2822 424866 -2586
rect 425102 -2822 444546 -2586
rect 444782 -2822 444866 -2586
rect 445102 -2822 464546 -2586
rect 464782 -2822 464866 -2586
rect 465102 -2822 484546 -2586
rect 484782 -2822 484866 -2586
rect 485102 -2822 504546 -2586
rect 504782 -2822 504866 -2586
rect 505102 -2822 524546 -2586
rect 524782 -2822 524866 -2586
rect 525102 -2822 544546 -2586
rect 544782 -2822 544866 -2586
rect 545102 -2822 564546 -2586
rect 564782 -2822 564866 -2586
rect 565102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 14546 -3226
rect 14782 -3462 14866 -3226
rect 15102 -3462 34546 -3226
rect 34782 -3462 34866 -3226
rect 35102 -3462 54546 -3226
rect 54782 -3462 54866 -3226
rect 55102 -3462 74546 -3226
rect 74782 -3462 74866 -3226
rect 75102 -3462 94546 -3226
rect 94782 -3462 94866 -3226
rect 95102 -3462 114546 -3226
rect 114782 -3462 114866 -3226
rect 115102 -3462 134546 -3226
rect 134782 -3462 134866 -3226
rect 135102 -3462 154546 -3226
rect 154782 -3462 154866 -3226
rect 155102 -3462 174546 -3226
rect 174782 -3462 174866 -3226
rect 175102 -3462 194546 -3226
rect 194782 -3462 194866 -3226
rect 195102 -3462 214546 -3226
rect 214782 -3462 214866 -3226
rect 215102 -3462 234546 -3226
rect 234782 -3462 234866 -3226
rect 235102 -3462 254546 -3226
rect 254782 -3462 254866 -3226
rect 255102 -3462 274546 -3226
rect 274782 -3462 274866 -3226
rect 275102 -3462 294546 -3226
rect 294782 -3462 294866 -3226
rect 295102 -3462 314546 -3226
rect 314782 -3462 314866 -3226
rect 315102 -3462 334546 -3226
rect 334782 -3462 334866 -3226
rect 335102 -3462 354546 -3226
rect 354782 -3462 354866 -3226
rect 355102 -3462 374546 -3226
rect 374782 -3462 374866 -3226
rect 375102 -3462 394546 -3226
rect 394782 -3462 394866 -3226
rect 395102 -3462 414546 -3226
rect 414782 -3462 414866 -3226
rect 415102 -3462 434546 -3226
rect 434782 -3462 434866 -3226
rect 435102 -3462 454546 -3226
rect 454782 -3462 454866 -3226
rect 455102 -3462 474546 -3226
rect 474782 -3462 474866 -3226
rect 475102 -3462 494546 -3226
rect 494782 -3462 494866 -3226
rect 495102 -3462 514546 -3226
rect 514782 -3462 514866 -3226
rect 515102 -3462 534546 -3226
rect 534782 -3462 534866 -3226
rect 535102 -3462 554546 -3226
rect 554782 -3462 554866 -3226
rect 555102 -3462 574546 -3226
rect 574782 -3462 574866 -3226
rect 575102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 14546 -3546
rect 14782 -3782 14866 -3546
rect 15102 -3782 34546 -3546
rect 34782 -3782 34866 -3546
rect 35102 -3782 54546 -3546
rect 54782 -3782 54866 -3546
rect 55102 -3782 74546 -3546
rect 74782 -3782 74866 -3546
rect 75102 -3782 94546 -3546
rect 94782 -3782 94866 -3546
rect 95102 -3782 114546 -3546
rect 114782 -3782 114866 -3546
rect 115102 -3782 134546 -3546
rect 134782 -3782 134866 -3546
rect 135102 -3782 154546 -3546
rect 154782 -3782 154866 -3546
rect 155102 -3782 174546 -3546
rect 174782 -3782 174866 -3546
rect 175102 -3782 194546 -3546
rect 194782 -3782 194866 -3546
rect 195102 -3782 214546 -3546
rect 214782 -3782 214866 -3546
rect 215102 -3782 234546 -3546
rect 234782 -3782 234866 -3546
rect 235102 -3782 254546 -3546
rect 254782 -3782 254866 -3546
rect 255102 -3782 274546 -3546
rect 274782 -3782 274866 -3546
rect 275102 -3782 294546 -3546
rect 294782 -3782 294866 -3546
rect 295102 -3782 314546 -3546
rect 314782 -3782 314866 -3546
rect 315102 -3782 334546 -3546
rect 334782 -3782 334866 -3546
rect 335102 -3782 354546 -3546
rect 354782 -3782 354866 -3546
rect 355102 -3782 374546 -3546
rect 374782 -3782 374866 -3546
rect 375102 -3782 394546 -3546
rect 394782 -3782 394866 -3546
rect 395102 -3782 414546 -3546
rect 414782 -3782 414866 -3546
rect 415102 -3782 434546 -3546
rect 434782 -3782 434866 -3546
rect 435102 -3782 454546 -3546
rect 454782 -3782 454866 -3546
rect 455102 -3782 474546 -3546
rect 474782 -3782 474866 -3546
rect 475102 -3782 494546 -3546
rect 494782 -3782 494866 -3546
rect 495102 -3782 514546 -3546
rect 514782 -3782 514866 -3546
rect 515102 -3782 534546 -3546
rect 534782 -3782 534866 -3546
rect 535102 -3782 554546 -3546
rect 554782 -3782 554866 -3546
rect 555102 -3782 574546 -3546
rect 574782 -3782 574866 -3546
rect 575102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 8266 -4186
rect 8502 -4422 8586 -4186
rect 8822 -4422 28266 -4186
rect 28502 -4422 28586 -4186
rect 28822 -4422 48266 -4186
rect 48502 -4422 48586 -4186
rect 48822 -4422 68266 -4186
rect 68502 -4422 68586 -4186
rect 68822 -4422 88266 -4186
rect 88502 -4422 88586 -4186
rect 88822 -4422 108266 -4186
rect 108502 -4422 108586 -4186
rect 108822 -4422 128266 -4186
rect 128502 -4422 128586 -4186
rect 128822 -4422 148266 -4186
rect 148502 -4422 148586 -4186
rect 148822 -4422 168266 -4186
rect 168502 -4422 168586 -4186
rect 168822 -4422 188266 -4186
rect 188502 -4422 188586 -4186
rect 188822 -4422 208266 -4186
rect 208502 -4422 208586 -4186
rect 208822 -4422 228266 -4186
rect 228502 -4422 228586 -4186
rect 228822 -4422 248266 -4186
rect 248502 -4422 248586 -4186
rect 248822 -4422 268266 -4186
rect 268502 -4422 268586 -4186
rect 268822 -4422 288266 -4186
rect 288502 -4422 288586 -4186
rect 288822 -4422 308266 -4186
rect 308502 -4422 308586 -4186
rect 308822 -4422 328266 -4186
rect 328502 -4422 328586 -4186
rect 328822 -4422 348266 -4186
rect 348502 -4422 348586 -4186
rect 348822 -4422 368266 -4186
rect 368502 -4422 368586 -4186
rect 368822 -4422 388266 -4186
rect 388502 -4422 388586 -4186
rect 388822 -4422 408266 -4186
rect 408502 -4422 408586 -4186
rect 408822 -4422 428266 -4186
rect 428502 -4422 428586 -4186
rect 428822 -4422 448266 -4186
rect 448502 -4422 448586 -4186
rect 448822 -4422 468266 -4186
rect 468502 -4422 468586 -4186
rect 468822 -4422 488266 -4186
rect 488502 -4422 488586 -4186
rect 488822 -4422 508266 -4186
rect 508502 -4422 508586 -4186
rect 508822 -4422 528266 -4186
rect 528502 -4422 528586 -4186
rect 528822 -4422 548266 -4186
rect 548502 -4422 548586 -4186
rect 548822 -4422 568266 -4186
rect 568502 -4422 568586 -4186
rect 568822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 8266 -4506
rect 8502 -4742 8586 -4506
rect 8822 -4742 28266 -4506
rect 28502 -4742 28586 -4506
rect 28822 -4742 48266 -4506
rect 48502 -4742 48586 -4506
rect 48822 -4742 68266 -4506
rect 68502 -4742 68586 -4506
rect 68822 -4742 88266 -4506
rect 88502 -4742 88586 -4506
rect 88822 -4742 108266 -4506
rect 108502 -4742 108586 -4506
rect 108822 -4742 128266 -4506
rect 128502 -4742 128586 -4506
rect 128822 -4742 148266 -4506
rect 148502 -4742 148586 -4506
rect 148822 -4742 168266 -4506
rect 168502 -4742 168586 -4506
rect 168822 -4742 188266 -4506
rect 188502 -4742 188586 -4506
rect 188822 -4742 208266 -4506
rect 208502 -4742 208586 -4506
rect 208822 -4742 228266 -4506
rect 228502 -4742 228586 -4506
rect 228822 -4742 248266 -4506
rect 248502 -4742 248586 -4506
rect 248822 -4742 268266 -4506
rect 268502 -4742 268586 -4506
rect 268822 -4742 288266 -4506
rect 288502 -4742 288586 -4506
rect 288822 -4742 308266 -4506
rect 308502 -4742 308586 -4506
rect 308822 -4742 328266 -4506
rect 328502 -4742 328586 -4506
rect 328822 -4742 348266 -4506
rect 348502 -4742 348586 -4506
rect 348822 -4742 368266 -4506
rect 368502 -4742 368586 -4506
rect 368822 -4742 388266 -4506
rect 388502 -4742 388586 -4506
rect 388822 -4742 408266 -4506
rect 408502 -4742 408586 -4506
rect 408822 -4742 428266 -4506
rect 428502 -4742 428586 -4506
rect 428822 -4742 448266 -4506
rect 448502 -4742 448586 -4506
rect 448822 -4742 468266 -4506
rect 468502 -4742 468586 -4506
rect 468822 -4742 488266 -4506
rect 488502 -4742 488586 -4506
rect 488822 -4742 508266 -4506
rect 508502 -4742 508586 -4506
rect 508822 -4742 528266 -4506
rect 528502 -4742 528586 -4506
rect 528822 -4742 548266 -4506
rect 548502 -4742 548586 -4506
rect 548822 -4742 568266 -4506
rect 568502 -4742 568586 -4506
rect 568822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 18266 -5146
rect 18502 -5382 18586 -5146
rect 18822 -5382 38266 -5146
rect 38502 -5382 38586 -5146
rect 38822 -5382 58266 -5146
rect 58502 -5382 58586 -5146
rect 58822 -5382 78266 -5146
rect 78502 -5382 78586 -5146
rect 78822 -5382 98266 -5146
rect 98502 -5382 98586 -5146
rect 98822 -5382 118266 -5146
rect 118502 -5382 118586 -5146
rect 118822 -5382 138266 -5146
rect 138502 -5382 138586 -5146
rect 138822 -5382 158266 -5146
rect 158502 -5382 158586 -5146
rect 158822 -5382 178266 -5146
rect 178502 -5382 178586 -5146
rect 178822 -5382 198266 -5146
rect 198502 -5382 198586 -5146
rect 198822 -5382 218266 -5146
rect 218502 -5382 218586 -5146
rect 218822 -5382 238266 -5146
rect 238502 -5382 238586 -5146
rect 238822 -5382 258266 -5146
rect 258502 -5382 258586 -5146
rect 258822 -5382 278266 -5146
rect 278502 -5382 278586 -5146
rect 278822 -5382 298266 -5146
rect 298502 -5382 298586 -5146
rect 298822 -5382 318266 -5146
rect 318502 -5382 318586 -5146
rect 318822 -5382 338266 -5146
rect 338502 -5382 338586 -5146
rect 338822 -5382 358266 -5146
rect 358502 -5382 358586 -5146
rect 358822 -5382 378266 -5146
rect 378502 -5382 378586 -5146
rect 378822 -5382 398266 -5146
rect 398502 -5382 398586 -5146
rect 398822 -5382 418266 -5146
rect 418502 -5382 418586 -5146
rect 418822 -5382 438266 -5146
rect 438502 -5382 438586 -5146
rect 438822 -5382 458266 -5146
rect 458502 -5382 458586 -5146
rect 458822 -5382 478266 -5146
rect 478502 -5382 478586 -5146
rect 478822 -5382 498266 -5146
rect 498502 -5382 498586 -5146
rect 498822 -5382 518266 -5146
rect 518502 -5382 518586 -5146
rect 518822 -5382 538266 -5146
rect 538502 -5382 538586 -5146
rect 538822 -5382 558266 -5146
rect 558502 -5382 558586 -5146
rect 558822 -5382 578266 -5146
rect 578502 -5382 578586 -5146
rect 578822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 18266 -5466
rect 18502 -5702 18586 -5466
rect 18822 -5702 38266 -5466
rect 38502 -5702 38586 -5466
rect 38822 -5702 58266 -5466
rect 58502 -5702 58586 -5466
rect 58822 -5702 78266 -5466
rect 78502 -5702 78586 -5466
rect 78822 -5702 98266 -5466
rect 98502 -5702 98586 -5466
rect 98822 -5702 118266 -5466
rect 118502 -5702 118586 -5466
rect 118822 -5702 138266 -5466
rect 138502 -5702 138586 -5466
rect 138822 -5702 158266 -5466
rect 158502 -5702 158586 -5466
rect 158822 -5702 178266 -5466
rect 178502 -5702 178586 -5466
rect 178822 -5702 198266 -5466
rect 198502 -5702 198586 -5466
rect 198822 -5702 218266 -5466
rect 218502 -5702 218586 -5466
rect 218822 -5702 238266 -5466
rect 238502 -5702 238586 -5466
rect 238822 -5702 258266 -5466
rect 258502 -5702 258586 -5466
rect 258822 -5702 278266 -5466
rect 278502 -5702 278586 -5466
rect 278822 -5702 298266 -5466
rect 298502 -5702 298586 -5466
rect 298822 -5702 318266 -5466
rect 318502 -5702 318586 -5466
rect 318822 -5702 338266 -5466
rect 338502 -5702 338586 -5466
rect 338822 -5702 358266 -5466
rect 358502 -5702 358586 -5466
rect 358822 -5702 378266 -5466
rect 378502 -5702 378586 -5466
rect 378822 -5702 398266 -5466
rect 398502 -5702 398586 -5466
rect 398822 -5702 418266 -5466
rect 418502 -5702 418586 -5466
rect 418822 -5702 438266 -5466
rect 438502 -5702 438586 -5466
rect 438822 -5702 458266 -5466
rect 458502 -5702 458586 -5466
rect 458822 -5702 478266 -5466
rect 478502 -5702 478586 -5466
rect 478822 -5702 498266 -5466
rect 498502 -5702 498586 -5466
rect 498822 -5702 518266 -5466
rect 518502 -5702 518586 -5466
rect 518822 -5702 538266 -5466
rect 538502 -5702 538586 -5466
rect 538822 -5702 558266 -5466
rect 558502 -5702 558586 -5466
rect 558822 -5702 578266 -5466
rect 578502 -5702 578586 -5466
rect 578822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 11986 -6106
rect 12222 -6342 12306 -6106
rect 12542 -6342 31986 -6106
rect 32222 -6342 32306 -6106
rect 32542 -6342 51986 -6106
rect 52222 -6342 52306 -6106
rect 52542 -6342 71986 -6106
rect 72222 -6342 72306 -6106
rect 72542 -6342 91986 -6106
rect 92222 -6342 92306 -6106
rect 92542 -6342 111986 -6106
rect 112222 -6342 112306 -6106
rect 112542 -6342 131986 -6106
rect 132222 -6342 132306 -6106
rect 132542 -6342 151986 -6106
rect 152222 -6342 152306 -6106
rect 152542 -6342 171986 -6106
rect 172222 -6342 172306 -6106
rect 172542 -6342 191986 -6106
rect 192222 -6342 192306 -6106
rect 192542 -6342 211986 -6106
rect 212222 -6342 212306 -6106
rect 212542 -6342 231986 -6106
rect 232222 -6342 232306 -6106
rect 232542 -6342 251986 -6106
rect 252222 -6342 252306 -6106
rect 252542 -6342 271986 -6106
rect 272222 -6342 272306 -6106
rect 272542 -6342 291986 -6106
rect 292222 -6342 292306 -6106
rect 292542 -6342 311986 -6106
rect 312222 -6342 312306 -6106
rect 312542 -6342 331986 -6106
rect 332222 -6342 332306 -6106
rect 332542 -6342 351986 -6106
rect 352222 -6342 352306 -6106
rect 352542 -6342 371986 -6106
rect 372222 -6342 372306 -6106
rect 372542 -6342 391986 -6106
rect 392222 -6342 392306 -6106
rect 392542 -6342 411986 -6106
rect 412222 -6342 412306 -6106
rect 412542 -6342 431986 -6106
rect 432222 -6342 432306 -6106
rect 432542 -6342 451986 -6106
rect 452222 -6342 452306 -6106
rect 452542 -6342 471986 -6106
rect 472222 -6342 472306 -6106
rect 472542 -6342 491986 -6106
rect 492222 -6342 492306 -6106
rect 492542 -6342 511986 -6106
rect 512222 -6342 512306 -6106
rect 512542 -6342 531986 -6106
rect 532222 -6342 532306 -6106
rect 532542 -6342 551986 -6106
rect 552222 -6342 552306 -6106
rect 552542 -6342 571986 -6106
rect 572222 -6342 572306 -6106
rect 572542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 11986 -6426
rect 12222 -6662 12306 -6426
rect 12542 -6662 31986 -6426
rect 32222 -6662 32306 -6426
rect 32542 -6662 51986 -6426
rect 52222 -6662 52306 -6426
rect 52542 -6662 71986 -6426
rect 72222 -6662 72306 -6426
rect 72542 -6662 91986 -6426
rect 92222 -6662 92306 -6426
rect 92542 -6662 111986 -6426
rect 112222 -6662 112306 -6426
rect 112542 -6662 131986 -6426
rect 132222 -6662 132306 -6426
rect 132542 -6662 151986 -6426
rect 152222 -6662 152306 -6426
rect 152542 -6662 171986 -6426
rect 172222 -6662 172306 -6426
rect 172542 -6662 191986 -6426
rect 192222 -6662 192306 -6426
rect 192542 -6662 211986 -6426
rect 212222 -6662 212306 -6426
rect 212542 -6662 231986 -6426
rect 232222 -6662 232306 -6426
rect 232542 -6662 251986 -6426
rect 252222 -6662 252306 -6426
rect 252542 -6662 271986 -6426
rect 272222 -6662 272306 -6426
rect 272542 -6662 291986 -6426
rect 292222 -6662 292306 -6426
rect 292542 -6662 311986 -6426
rect 312222 -6662 312306 -6426
rect 312542 -6662 331986 -6426
rect 332222 -6662 332306 -6426
rect 332542 -6662 351986 -6426
rect 352222 -6662 352306 -6426
rect 352542 -6662 371986 -6426
rect 372222 -6662 372306 -6426
rect 372542 -6662 391986 -6426
rect 392222 -6662 392306 -6426
rect 392542 -6662 411986 -6426
rect 412222 -6662 412306 -6426
rect 412542 -6662 431986 -6426
rect 432222 -6662 432306 -6426
rect 432542 -6662 451986 -6426
rect 452222 -6662 452306 -6426
rect 452542 -6662 471986 -6426
rect 472222 -6662 472306 -6426
rect 472542 -6662 491986 -6426
rect 492222 -6662 492306 -6426
rect 492542 -6662 511986 -6426
rect 512222 -6662 512306 -6426
rect 512542 -6662 531986 -6426
rect 532222 -6662 532306 -6426
rect 532542 -6662 551986 -6426
rect 552222 -6662 552306 -6426
rect 552542 -6662 571986 -6426
rect 572222 -6662 572306 -6426
rect 572542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 21986 -7066
rect 22222 -7302 22306 -7066
rect 22542 -7302 41986 -7066
rect 42222 -7302 42306 -7066
rect 42542 -7302 61986 -7066
rect 62222 -7302 62306 -7066
rect 62542 -7302 81986 -7066
rect 82222 -7302 82306 -7066
rect 82542 -7302 101986 -7066
rect 102222 -7302 102306 -7066
rect 102542 -7302 121986 -7066
rect 122222 -7302 122306 -7066
rect 122542 -7302 141986 -7066
rect 142222 -7302 142306 -7066
rect 142542 -7302 161986 -7066
rect 162222 -7302 162306 -7066
rect 162542 -7302 181986 -7066
rect 182222 -7302 182306 -7066
rect 182542 -7302 201986 -7066
rect 202222 -7302 202306 -7066
rect 202542 -7302 221986 -7066
rect 222222 -7302 222306 -7066
rect 222542 -7302 241986 -7066
rect 242222 -7302 242306 -7066
rect 242542 -7302 261986 -7066
rect 262222 -7302 262306 -7066
rect 262542 -7302 281986 -7066
rect 282222 -7302 282306 -7066
rect 282542 -7302 301986 -7066
rect 302222 -7302 302306 -7066
rect 302542 -7302 321986 -7066
rect 322222 -7302 322306 -7066
rect 322542 -7302 341986 -7066
rect 342222 -7302 342306 -7066
rect 342542 -7302 361986 -7066
rect 362222 -7302 362306 -7066
rect 362542 -7302 381986 -7066
rect 382222 -7302 382306 -7066
rect 382542 -7302 401986 -7066
rect 402222 -7302 402306 -7066
rect 402542 -7302 421986 -7066
rect 422222 -7302 422306 -7066
rect 422542 -7302 441986 -7066
rect 442222 -7302 442306 -7066
rect 442542 -7302 461986 -7066
rect 462222 -7302 462306 -7066
rect 462542 -7302 481986 -7066
rect 482222 -7302 482306 -7066
rect 482542 -7302 501986 -7066
rect 502222 -7302 502306 -7066
rect 502542 -7302 521986 -7066
rect 522222 -7302 522306 -7066
rect 522542 -7302 541986 -7066
rect 542222 -7302 542306 -7066
rect 542542 -7302 561986 -7066
rect 562222 -7302 562306 -7066
rect 562542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 21986 -7386
rect 22222 -7622 22306 -7386
rect 22542 -7622 41986 -7386
rect 42222 -7622 42306 -7386
rect 42542 -7622 61986 -7386
rect 62222 -7622 62306 -7386
rect 62542 -7622 81986 -7386
rect 82222 -7622 82306 -7386
rect 82542 -7622 101986 -7386
rect 102222 -7622 102306 -7386
rect 102542 -7622 121986 -7386
rect 122222 -7622 122306 -7386
rect 122542 -7622 141986 -7386
rect 142222 -7622 142306 -7386
rect 142542 -7622 161986 -7386
rect 162222 -7622 162306 -7386
rect 162542 -7622 181986 -7386
rect 182222 -7622 182306 -7386
rect 182542 -7622 201986 -7386
rect 202222 -7622 202306 -7386
rect 202542 -7622 221986 -7386
rect 222222 -7622 222306 -7386
rect 222542 -7622 241986 -7386
rect 242222 -7622 242306 -7386
rect 242542 -7622 261986 -7386
rect 262222 -7622 262306 -7386
rect 262542 -7622 281986 -7386
rect 282222 -7622 282306 -7386
rect 282542 -7622 301986 -7386
rect 302222 -7622 302306 -7386
rect 302542 -7622 321986 -7386
rect 322222 -7622 322306 -7386
rect 322542 -7622 341986 -7386
rect 342222 -7622 342306 -7386
rect 342542 -7622 361986 -7386
rect 362222 -7622 362306 -7386
rect 362542 -7622 381986 -7386
rect 382222 -7622 382306 -7386
rect 382542 -7622 401986 -7386
rect 402222 -7622 402306 -7386
rect 402542 -7622 421986 -7386
rect 422222 -7622 422306 -7386
rect 422542 -7622 441986 -7386
rect 442222 -7622 442306 -7386
rect 442542 -7622 461986 -7386
rect 462222 -7622 462306 -7386
rect 462542 -7622 481986 -7386
rect 482222 -7622 482306 -7386
rect 482542 -7622 501986 -7386
rect 502222 -7622 502306 -7386
rect 502542 -7622 521986 -7386
rect 522222 -7622 522306 -7386
rect 522542 -7622 541986 -7386
rect 542222 -7622 542306 -7386
rect 542542 -7622 561986 -7386
rect 562222 -7622 562306 -7386
rect 562542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use to_ALU_opt_TMR_KP_Voter  TMR_ALU
timestamp 1640855983
transform 1 0 20000 0 1 20000
box 0 0 50151 52295
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 20794 -1894 21414 18000 6 vccd1
port 531 nsew power input
rlabel metal4 s 40794 -1894 41414 18000 6 vccd1
port 531 nsew power input
rlabel metal4 s 60794 -1894 61414 18000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 794 -1894 1414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 20794 74295 21414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 40794 74295 41414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 60794 74295 61414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 80794 -1894 81414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 100794 -1894 101414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 120794 -1894 121414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 140794 -1894 141414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 160794 -1894 161414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 180794 -1894 181414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 200794 -1894 201414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 220794 -1894 221414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 240794 -1894 241414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 260794 -1894 261414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 280794 -1894 281414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 300794 -1894 301414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 320794 -1894 321414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 340794 -1894 341414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 360794 -1894 361414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 380794 -1894 381414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 400794 -1894 401414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 420794 -1894 421414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 440794 -1894 441414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 460794 -1894 461414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 480794 -1894 481414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 500794 -1894 501414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 520794 -1894 521414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 540794 -1894 541414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 560794 -1894 561414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 580794 -1894 581414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 24514 -3814 25134 18000 6 vccd2
port 532 nsew power input
rlabel metal4 s 44514 -3814 45134 18000 6 vccd2
port 532 nsew power input
rlabel metal4 s 64514 -3814 65134 18000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 4514 -3814 5134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 24514 74295 25134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 44514 74295 45134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 64514 74295 65134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 84514 -3814 85134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 104514 -3814 105134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 124514 -3814 125134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 144514 -3814 145134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 164514 -3814 165134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 184514 -3814 185134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 204514 -3814 205134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 224514 -3814 225134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 244514 -3814 245134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 264514 -3814 265134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 284514 -3814 285134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 304514 -3814 305134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 324514 -3814 325134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 344514 -3814 345134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 364514 -3814 365134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 384514 -3814 385134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 404514 -3814 405134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 424514 -3814 425134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 444514 -3814 445134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 464514 -3814 465134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 484514 -3814 485134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 504514 -3814 505134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 524514 -3814 525134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 544514 -3814 545134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 564514 -3814 565134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 28234 -5734 28854 18000 6 vdda1
port 533 nsew power input
rlabel metal4 s 48234 -5734 48854 18000 6 vdda1
port 533 nsew power input
rlabel metal4 s 68234 -5734 68854 18000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 8234 -5734 8854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 28234 74295 28854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 48234 74295 48854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 68234 74295 68854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 88234 -5734 88854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 108234 -5734 108854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 128234 -5734 128854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 148234 -5734 148854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 168234 -5734 168854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 188234 -5734 188854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 208234 -5734 208854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 228234 -5734 228854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 248234 -5734 248854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 268234 -5734 268854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 288234 -5734 288854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 308234 -5734 308854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 328234 -5734 328854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 348234 -5734 348854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 368234 -5734 368854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 388234 -5734 388854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 408234 -5734 408854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 428234 -5734 428854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 448234 -5734 448854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 468234 -5734 468854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 488234 -5734 488854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 508234 -5734 508854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 528234 -5734 528854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 548234 -5734 548854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 568234 -5734 568854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 31954 -7654 32574 18000 6 vdda2
port 534 nsew power input
rlabel metal4 s 51954 -7654 52574 18000 6 vdda2
port 534 nsew power input
rlabel metal4 s 71954 -7654 72574 18000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 11954 -7654 12574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 31954 74295 32574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 51954 74295 52574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 71954 74295 72574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 91954 -7654 92574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 111954 -7654 112574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 131954 -7654 132574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 151954 -7654 152574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 171954 -7654 172574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 191954 -7654 192574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 211954 -7654 212574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 231954 -7654 232574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 251954 -7654 252574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 271954 -7654 272574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 291954 -7654 292574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 311954 -7654 312574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 331954 -7654 332574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 351954 -7654 352574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 371954 -7654 372574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 391954 -7654 392574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 411954 -7654 412574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 431954 -7654 432574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 451954 -7654 452574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 471954 -7654 472574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 491954 -7654 492574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 511954 -7654 512574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 531954 -7654 532574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 551954 -7654 552574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 571954 -7654 572574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 18234 -5734 18854 18000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 38234 -5734 38854 18000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 58234 -5734 58854 18000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 18234 74295 18854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 38234 74295 38854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 58234 74295 58854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 78234 -5734 78854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98234 -5734 98854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 118234 -5734 118854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 138234 -5734 138854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 158234 -5734 158854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 178234 -5734 178854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 198234 -5734 198854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 218234 -5734 218854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 238234 -5734 238854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 258234 -5734 258854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 278234 -5734 278854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 298234 -5734 298854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 318234 -5734 318854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 338234 -5734 338854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 358234 -5734 358854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 378234 -5734 378854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 398234 -5734 398854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 418234 -5734 418854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 438234 -5734 438854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 458234 -5734 458854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 478234 -5734 478854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 498234 -5734 498854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 518234 -5734 518854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 538234 -5734 538854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 558234 -5734 558854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 578234 -5734 578854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 21954 -7654 22574 18000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 41954 -7654 42574 18000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 61954 -7654 62574 18000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 21954 74295 22574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 41954 74295 42574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 61954 74295 62574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 81954 -7654 82574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101954 -7654 102574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 121954 -7654 122574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 141954 -7654 142574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 161954 -7654 162574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 181954 -7654 182574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 201954 -7654 202574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 221954 -7654 222574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 241954 -7654 242574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 261954 -7654 262574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 281954 -7654 282574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 301954 -7654 302574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 321954 -7654 322574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 341954 -7654 342574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 361954 -7654 362574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 381954 -7654 382574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 401954 -7654 402574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 421954 -7654 422574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 441954 -7654 442574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 461954 -7654 462574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 481954 -7654 482574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 501954 -7654 502574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 521954 -7654 522574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 541954 -7654 542574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 561954 -7654 562574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 30794 -1894 31414 18000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 50794 -1894 51414 18000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 70794 -1894 71414 18000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 10794 -1894 11414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 30794 74295 31414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 50794 74295 51414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 70794 74295 71414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90794 -1894 91414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 110794 -1894 111414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 130794 -1894 131414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 150794 -1894 151414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 170794 -1894 171414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 190794 -1894 191414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 210794 -1894 211414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 230794 -1894 231414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 250794 -1894 251414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 270794 -1894 271414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 290794 -1894 291414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 310794 -1894 311414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 330794 -1894 331414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 350794 -1894 351414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 370794 -1894 371414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 390794 -1894 391414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 410794 -1894 411414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 430794 -1894 431414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 450794 -1894 451414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 470794 -1894 471414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 490794 -1894 491414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 510794 -1894 511414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 530794 -1894 531414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 550794 -1894 551414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 570794 -1894 571414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 34514 -3814 35134 18000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 54514 -3814 55134 18000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 14514 -3814 15134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 34514 74295 35134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 54514 74295 55134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 74514 -3814 75134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94514 -3814 95134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 114514 -3814 115134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 134514 -3814 135134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 154514 -3814 155134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 174514 -3814 175134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 194514 -3814 195134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 214514 -3814 215134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 234514 -3814 235134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 254514 -3814 255134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 274514 -3814 275134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 294514 -3814 295134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 314514 -3814 315134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 334514 -3814 335134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 354514 -3814 355134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 374514 -3814 375134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 394514 -3814 395134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 414514 -3814 415134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 434514 -3814 435134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 454514 -3814 455134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 474514 -3814 475134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 494514 -3814 495134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 514514 -3814 515134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 534514 -3814 535134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 554514 -3814 555134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 574514 -3814 575134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
